module tb ();
   
   logic[23:0]  N, D;
   logic[23:0]  Out;
   logic[2:0]   Ma, Mb;
   logic        Sn, Sd, Ms, Mq, La, Lb, Lk, Lf, clk;
   
  // instantiate device under test
  main dut (N, D, Sn, Sd, Mb, Ma, Ms, Mq, La, Lb, Lk, Lf, clk, Out);

  /*/ generate clock
  always 
    begin
      clk = 1; #10; clk = 0; #10;
    end
  */  
   integer STest, errorCount;
   initial
     begin
        $display ("Testing... ");
        
        #0 errorCount = 0;
		#0 Lf = 1'b0;
        
        //Cycle 0
        #0  N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
		#0  clk = 1;
        #10  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
		#0  clk = 0;
		#10
	
        //Cycle 1
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
		#0  clk = 1;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
		#10
        
        //Cycle 2
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
		#0  clk = 1;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 3
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
       
        
        //Cycle 4
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 5
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 6
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 7
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 8
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 9
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 10
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 11
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Final
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        assert (Out == 24'b110000000000000000000000) else begin
            $error ("Crap");
            end
        
        //Cycle 0
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10

		
        //Cycle 1
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 2
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 3
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
       
        
        //Cycle 4
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        
        //Cycle 5
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 6
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        
        //Cycle 7
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 8
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 9
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 10
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 11
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Final
        #0 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        assert (Out == 24'b100000000000000000000000) else begin
            $error ("Crap Again");
            end
        
        //Cycle 0
        #0 N = 24'b111100000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10

        //Cycle 1
        #0 N = 24'b111100000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 3'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 2
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 3
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
       
        
        //Cycle 4
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 5
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 6
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 7
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 8
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 9
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 10
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 11
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Final
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        assert (Out == 24'b101000000000000000000000) else begin
            $error ("Crap x3");
            end
			
		//Inverse of test 3
		//Cycle 0
		#0 Lf = 1'b1;
		#0 clk = 1;
		#10 Lf = 1'b0;
		#0 clk = 0;
		
        #0  Mb = 3'd3;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10

        //Cycle 1
        #0  Mb = 3'd0;
        #0  Ma = 3'd6;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 2
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 3
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
		#0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
       
        
        //Cycle 4
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 5
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 6
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 7
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 8
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 9
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 10
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 11
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Final
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        assert (Out == 24'b011001100110011001100110) else begin
            $error ("Crap x3 - Inverse");
            end
		
        
         
        //Cycle 0
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd0;
        #0  Ma = 3'd5;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10

        //Cycle 1
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd0;
        #0  Ma = 3'd0;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 2
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd0;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 3
        #0  N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 4
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 5
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 6
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 7
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 8
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 9
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 10
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Cycle 11
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 12
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 13
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 14
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 15
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 16
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
		
        //Cycle 17
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        //Final
        #0 N = 24'b110000000000000000000000;
        #0  Mb = 3'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 1;
		#10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #0  clk = 0;
        #10
        
        assert (Out == 24'b100111001100010001110000) else begin
            $error ("Crap x4");
            end
        
    end
        
endmodule
