module tb ();
   
   logic[23:0]  N, D;
   logic[26:0]  Out;
   logic[2:0]   Ma;
   logic[1:0]   Mb;
   logic        Sn, Sd, Ms, Mq, La, Lb, Lk, clk;
   
  // instantiate device under test
  main dut (N, D, Sn, Sd, Mb, Ma, Ms, Mq, La, Lb, Lk, clk, Out);

  // generate clock
  always 
    begin
      clk = 1; #10; clk = 0; #10;
    end
    
   integer STest, errorCount;
   initial
     begin
        $display ("Testing... ");
        
        errorCount = 0;
        
        //Cycle 0
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        //STest = 27'b000000000000;
        //assert (Out == STest) else begin 
          //  $error("ERROR! Value N = %0d, D = %0d, \nS:%0d  !=  STest: %0d\n", N, D, Out, STest);
           // errorCount++;
            //end
        //Cycle 1
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #10  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 2
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #10  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #15  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 3
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
       
        
        //Cycle 4
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 5
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 6
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 7
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 8
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 9
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 10
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 11
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Final
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        assert (Out == 24'b110000000000000000000000) else begin
            $error ("Crap");
            end
        #10 
        //Cycle 0
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        //STest = 27'b000000000000;
        //assert (Out == STest) else begin 
          //  $error("ERROR! Value N = %0d, D = %0d, \nS:%0d  !=  STest: %0d\n", N, D, Out, STest);
           // errorCount++;
            //end
        //Cycle 1
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #10  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 2
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #10  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #15  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 3
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
       
        
        //Cycle 4
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 5
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 6
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 7
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 8
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 9
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 10
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 11
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Final
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        assert (Out == 24'b100000000000000000000000) else begin
            $error ("Crap Again");
            end
            
        #10 
        //Cycle 0
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd1;
        #0  Ma = 3'd5;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5

        //Cycle 1
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd0;
        #0  Ma = 3'd1;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #5  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #10  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 2
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #10  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #15  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 3
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
       
        
        //Cycle 4
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 5
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 6
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 7
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 8
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 9
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 10
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 11
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Final
        #20 N = 24'b110000000000000000000000;
        #0  D = 24'b100110011001100110011001;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b0;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        assert (Out == 24'b101000000000000000000000) else begin
            $error ("Crap x3");
            end
        
        #10 
        //Cycle 0
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd0;
        #0  Ma = 3'd5;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #5  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        #10 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5

        //Cycle 1
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd0;
        #0  Ma = 3'd0;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #5  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #10  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 2
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd0;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #10 La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        #15 La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        #5
        
        //Cycle 3
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
       
        
        //Cycle 4
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 5
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 6
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        
        
        //Cycle 7
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 8
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b1;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Cycle 9
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        
        
        //Cycle 10
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        //Cycle 11
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        //Cycle 12
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        
        //Cycle 13
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        //Cycle 14
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        //Cycle 15
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b1;
        
        //Cycle 16
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd4;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b1;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        //Cycle 17
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd3;
        #0  Ms = 1'b1;
        #0  Mq = 1'b0;
        #0  La = 1'b0;
        #0  Lb = 1'b1;
        #0  Lk = 1'b1;
        
        
        //Final
        #20 N = 24'b110000000000000000000000;
        #0  Mb = 2'd2;
        #0  Ma = 3'd2;
        #0  Ms = 1'b1;
        #0  Mq = 1'b1;
        #0  La = 1'b0;
        #0  Lb = 1'b0;
        #0  Lk = 1'b0;
        
        
        assert (Out == 24'b100111001100010001110000) else begin
            $error ("Crap x4");
            end
        
    end
        
endmodule
