module multiplier (Z, X, Y);
	
	input logic [26:0] Y;
	input logic [26:0] X;
	output logic [53:0] Z;


	logic [26:0] P0;
	logic [26:0] carry1;
	logic [26:0] sum1;
	logic [26:0] P1;
	logic [26:0] carry2;
	logic [26:0] sum2;
	logic [26:0] P2;
	logic [26:0] carry3;
	logic [26:0] sum3;
	logic [26:0] P3;
	logic [26:0] carry4;
	logic [26:0] sum4;
	logic [26:0] P4;
	logic [26:0] carry5;
	logic [26:0] sum5;
	logic [26:0] P5;
	logic [26:0] carry6;
	logic [26:0] sum6;
	logic [26:0] P6;
	logic [26:0] carry7;
	logic [26:0] sum7;
	logic [26:0] P7;
	logic [26:0] carry8;
	logic [26:0] sum8;
	logic [26:0] P8;
	logic [26:0] carry9;
	logic [26:0] sum9;
	logic [26:0] P9;
	logic [26:0] carry10;
	logic [26:0] sum10;
	logic [26:0] P10;
	logic [26:0] carry11;
	logic [26:0] sum11;
	logic [26:0] P11;
	logic [26:0] carry12;
	logic [26:0] sum12;
	logic [26:0] P12;
	logic [26:0] carry13;
	logic [26:0] sum13;
	logic [26:0] P13;
	logic [26:0] carry14;
	logic [26:0] sum14;
	logic [26:0] P14;
	logic [26:0] carry15;
	logic [26:0] sum15;
	logic [26:0] P15;
	logic [26:0] carry16;
	logic [26:0] sum16;
	logic [26:0] P16;
	logic [26:0] carry17;
	logic [26:0] sum17;
	logic [26:0] P17;
	logic [26:0] carry18;
	logic [26:0] sum18;
	logic [26:0] P18;
	logic [26:0] carry19;
	logic [26:0] sum19;
	logic [26:0] P19;
	logic [26:0] carry20;
	logic [26:0] sum20;
	logic [26:0] P20;
	logic [26:0] carry21;
	logic [26:0] sum21;
	logic [26:0] P21;
	logic [26:0] carry22;
	logic [26:0] sum22;
	logic [26:0] P22;
	logic [26:0] carry23;
	logic [26:0] sum23;
	logic [26:0] P23;
	logic [26:0] carry24;
	logic [26:0] sum24;
	logic [26:0] P24;
	logic [26:0] carry25;
	logic [26:0] sum25;
	logic [26:0] P25;
	logic [26:0] carry26;
	logic [26:0] sum26;
	logic [26:0] P26;
	logic [26:0] carry27;
	logic [26:0] sum27;
	logic [52:0] carry28;


	// generate the partial products.
	and pp1(P0[26], X[26], Y[0]);
	and pp2(P0[25], X[25], Y[0]);
	and pp3(P0[24], X[24], Y[0]);
	and pp4(P0[23], X[23], Y[0]);
	and pp5(P0[22], X[22], Y[0]);
	and pp6(P0[21], X[21], Y[0]);
	and pp7(P0[20], X[20], Y[0]);
	and pp8(P0[19], X[19], Y[0]);
	and pp9(P0[18], X[18], Y[0]);
	and pp10(P0[17], X[17], Y[0]);
	and pp11(P0[16], X[16], Y[0]);
	and pp12(P0[15], X[15], Y[0]);
	and pp13(P0[14], X[14], Y[0]);
	and pp14(P0[13], X[13], Y[0]);
	and pp15(P0[12], X[12], Y[0]);
	and pp16(P0[11], X[11], Y[0]);
	and pp17(P0[10], X[10], Y[0]);
	and pp18(P0[9], X[9], Y[0]);
	and pp19(P0[8], X[8], Y[0]);
	and pp20(P0[7], X[7], Y[0]);
	and pp21(P0[6], X[6], Y[0]);
	and pp22(P0[5], X[5], Y[0]);
	and pp23(P0[4], X[4], Y[0]);
	and pp24(P0[3], X[3], Y[0]);
	and pp25(P0[2], X[2], Y[0]);
	and pp26(P0[1], X[1], Y[0]);
	and pp27(P0[0], X[0], Y[0]);
	and pp28(sum1[26], X[26], Y[1]);
	and pp29(P1[25], X[25], Y[1]);
	and pp30(P1[24], X[24], Y[1]);
	and pp31(P1[23], X[23], Y[1]);
	and pp32(P1[22], X[22], Y[1]);
	and pp33(P1[21], X[21], Y[1]);
	and pp34(P1[20], X[20], Y[1]);
	and pp35(P1[19], X[19], Y[1]);
	and pp36(P1[18], X[18], Y[1]);
	and pp37(P1[17], X[17], Y[1]);
	and pp38(P1[16], X[16], Y[1]);
	and pp39(P1[15], X[15], Y[1]);
	and pp40(P1[14], X[14], Y[1]);
	and pp41(P1[13], X[13], Y[1]);
	and pp42(P1[12], X[12], Y[1]);
	and pp43(P1[11], X[11], Y[1]);
	and pp44(P1[10], X[10], Y[1]);
	and pp45(P1[9], X[9], Y[1]);
	and pp46(P1[8], X[8], Y[1]);
	and pp47(P1[7], X[7], Y[1]);
	and pp48(P1[6], X[6], Y[1]);
	and pp49(P1[5], X[5], Y[1]);
	and pp50(P1[4], X[4], Y[1]);
	and pp51(P1[3], X[3], Y[1]);
	and pp52(P1[2], X[2], Y[1]);
	and pp53(P1[1], X[1], Y[1]);
	and pp54(P1[0], X[0], Y[1]);
	and pp55(sum2[26], X[26], Y[2]);
	and pp56(P2[25], X[25], Y[2]);
	and pp57(P2[24], X[24], Y[2]);
	and pp58(P2[23], X[23], Y[2]);
	and pp59(P2[22], X[22], Y[2]);
	and pp60(P2[21], X[21], Y[2]);
	and pp61(P2[20], X[20], Y[2]);
	and pp62(P2[19], X[19], Y[2]);
	and pp63(P2[18], X[18], Y[2]);
	and pp64(P2[17], X[17], Y[2]);
	and pp65(P2[16], X[16], Y[2]);
	and pp66(P2[15], X[15], Y[2]);
	and pp67(P2[14], X[14], Y[2]);
	and pp68(P2[13], X[13], Y[2]);
	and pp69(P2[12], X[12], Y[2]);
	and pp70(P2[11], X[11], Y[2]);
	and pp71(P2[10], X[10], Y[2]);
	and pp72(P2[9], X[9], Y[2]);
	and pp73(P2[8], X[8], Y[2]);
	and pp74(P2[7], X[7], Y[2]);
	and pp75(P2[6], X[6], Y[2]);
	and pp76(P2[5], X[5], Y[2]);
	and pp77(P2[4], X[4], Y[2]);
	and pp78(P2[3], X[3], Y[2]);
	and pp79(P2[2], X[2], Y[2]);
	and pp80(P2[1], X[1], Y[2]);
	and pp81(P2[0], X[0], Y[2]);
	and pp82(sum3[26], X[26], Y[3]);
	and pp83(P3[25], X[25], Y[3]);
	and pp84(P3[24], X[24], Y[3]);
	and pp85(P3[23], X[23], Y[3]);
	and pp86(P3[22], X[22], Y[3]);
	and pp87(P3[21], X[21], Y[3]);
	and pp88(P3[20], X[20], Y[3]);
	and pp89(P3[19], X[19], Y[3]);
	and pp90(P3[18], X[18], Y[3]);
	and pp91(P3[17], X[17], Y[3]);
	and pp92(P3[16], X[16], Y[3]);
	and pp93(P3[15], X[15], Y[3]);
	and pp94(P3[14], X[14], Y[3]);
	and pp95(P3[13], X[13], Y[3]);
	and pp96(P3[12], X[12], Y[3]);
	and pp97(P3[11], X[11], Y[3]);
	and pp98(P3[10], X[10], Y[3]);
	and pp99(P3[9], X[9], Y[3]);
	and pp100(P3[8], X[8], Y[3]);
	and pp101(P3[7], X[7], Y[3]);
	and pp102(P3[6], X[6], Y[3]);
	and pp103(P3[5], X[5], Y[3]);
	and pp104(P3[4], X[4], Y[3]);
	and pp105(P3[3], X[3], Y[3]);
	and pp106(P3[2], X[2], Y[3]);
	and pp107(P3[1], X[1], Y[3]);
	and pp108(P3[0], X[0], Y[3]);
	and pp109(sum4[26], X[26], Y[4]);
	and pp110(P4[25], X[25], Y[4]);
	and pp111(P4[24], X[24], Y[4]);
	and pp112(P4[23], X[23], Y[4]);
	and pp113(P4[22], X[22], Y[4]);
	and pp114(P4[21], X[21], Y[4]);
	and pp115(P4[20], X[20], Y[4]);
	and pp116(P4[19], X[19], Y[4]);
	and pp117(P4[18], X[18], Y[4]);
	and pp118(P4[17], X[17], Y[4]);
	and pp119(P4[16], X[16], Y[4]);
	and pp120(P4[15], X[15], Y[4]);
	and pp121(P4[14], X[14], Y[4]);
	and pp122(P4[13], X[13], Y[4]);
	and pp123(P4[12], X[12], Y[4]);
	and pp124(P4[11], X[11], Y[4]);
	and pp125(P4[10], X[10], Y[4]);
	and pp126(P4[9], X[9], Y[4]);
	and pp127(P4[8], X[8], Y[4]);
	and pp128(P4[7], X[7], Y[4]);
	and pp129(P4[6], X[6], Y[4]);
	and pp130(P4[5], X[5], Y[4]);
	and pp131(P4[4], X[4], Y[4]);
	and pp132(P4[3], X[3], Y[4]);
	and pp133(P4[2], X[2], Y[4]);
	and pp134(P4[1], X[1], Y[4]);
	and pp135(P4[0], X[0], Y[4]);
	and pp136(sum5[26], X[26], Y[5]);
	and pp137(P5[25], X[25], Y[5]);
	and pp138(P5[24], X[24], Y[5]);
	and pp139(P5[23], X[23], Y[5]);
	and pp140(P5[22], X[22], Y[5]);
	and pp141(P5[21], X[21], Y[5]);
	and pp142(P5[20], X[20], Y[5]);
	and pp143(P5[19], X[19], Y[5]);
	and pp144(P5[18], X[18], Y[5]);
	and pp145(P5[17], X[17], Y[5]);
	and pp146(P5[16], X[16], Y[5]);
	and pp147(P5[15], X[15], Y[5]);
	and pp148(P5[14], X[14], Y[5]);
	and pp149(P5[13], X[13], Y[5]);
	and pp150(P5[12], X[12], Y[5]);
	and pp151(P5[11], X[11], Y[5]);
	and pp152(P5[10], X[10], Y[5]);
	and pp153(P5[9], X[9], Y[5]);
	and pp154(P5[8], X[8], Y[5]);
	and pp155(P5[7], X[7], Y[5]);
	and pp156(P5[6], X[6], Y[5]);
	and pp157(P5[5], X[5], Y[5]);
	and pp158(P5[4], X[4], Y[5]);
	and pp159(P5[3], X[3], Y[5]);
	and pp160(P5[2], X[2], Y[5]);
	and pp161(P5[1], X[1], Y[5]);
	and pp162(P5[0], X[0], Y[5]);
	and pp163(sum6[26], X[26], Y[6]);
	and pp164(P6[25], X[25], Y[6]);
	and pp165(P6[24], X[24], Y[6]);
	and pp166(P6[23], X[23], Y[6]);
	and pp167(P6[22], X[22], Y[6]);
	and pp168(P6[21], X[21], Y[6]);
	and pp169(P6[20], X[20], Y[6]);
	and pp170(P6[19], X[19], Y[6]);
	and pp171(P6[18], X[18], Y[6]);
	and pp172(P6[17], X[17], Y[6]);
	and pp173(P6[16], X[16], Y[6]);
	and pp174(P6[15], X[15], Y[6]);
	and pp175(P6[14], X[14], Y[6]);
	and pp176(P6[13], X[13], Y[6]);
	and pp177(P6[12], X[12], Y[6]);
	and pp178(P6[11], X[11], Y[6]);
	and pp179(P6[10], X[10], Y[6]);
	and pp180(P6[9], X[9], Y[6]);
	and pp181(P6[8], X[8], Y[6]);
	and pp182(P6[7], X[7], Y[6]);
	and pp183(P6[6], X[6], Y[6]);
	and pp184(P6[5], X[5], Y[6]);
	and pp185(P6[4], X[4], Y[6]);
	and pp186(P6[3], X[3], Y[6]);
	and pp187(P6[2], X[2], Y[6]);
	and pp188(P6[1], X[1], Y[6]);
	and pp189(P6[0], X[0], Y[6]);
	and pp190(sum7[26], X[26], Y[7]);
	and pp191(P7[25], X[25], Y[7]);
	and pp192(P7[24], X[24], Y[7]);
	and pp193(P7[23], X[23], Y[7]);
	and pp194(P7[22], X[22], Y[7]);
	and pp195(P7[21], X[21], Y[7]);
	and pp196(P7[20], X[20], Y[7]);
	and pp197(P7[19], X[19], Y[7]);
	and pp198(P7[18], X[18], Y[7]);
	and pp199(P7[17], X[17], Y[7]);
	and pp200(P7[16], X[16], Y[7]);
	and pp201(P7[15], X[15], Y[7]);
	and pp202(P7[14], X[14], Y[7]);
	and pp203(P7[13], X[13], Y[7]);
	and pp204(P7[12], X[12], Y[7]);
	and pp205(P7[11], X[11], Y[7]);
	and pp206(P7[10], X[10], Y[7]);
	and pp207(P7[9], X[9], Y[7]);
	and pp208(P7[8], X[8], Y[7]);
	and pp209(P7[7], X[7], Y[7]);
	and pp210(P7[6], X[6], Y[7]);
	and pp211(P7[5], X[5], Y[7]);
	and pp212(P7[4], X[4], Y[7]);
	and pp213(P7[3], X[3], Y[7]);
	and pp214(P7[2], X[2], Y[7]);
	and pp215(P7[1], X[1], Y[7]);
	and pp216(P7[0], X[0], Y[7]);
	and pp217(sum8[26], X[26], Y[8]);
	and pp218(P8[25], X[25], Y[8]);
	and pp219(P8[24], X[24], Y[8]);
	and pp220(P8[23], X[23], Y[8]);
	and pp221(P8[22], X[22], Y[8]);
	and pp222(P8[21], X[21], Y[8]);
	and pp223(P8[20], X[20], Y[8]);
	and pp224(P8[19], X[19], Y[8]);
	and pp225(P8[18], X[18], Y[8]);
	and pp226(P8[17], X[17], Y[8]);
	and pp227(P8[16], X[16], Y[8]);
	and pp228(P8[15], X[15], Y[8]);
	and pp229(P8[14], X[14], Y[8]);
	and pp230(P8[13], X[13], Y[8]);
	and pp231(P8[12], X[12], Y[8]);
	and pp232(P8[11], X[11], Y[8]);
	and pp233(P8[10], X[10], Y[8]);
	and pp234(P8[9], X[9], Y[8]);
	and pp235(P8[8], X[8], Y[8]);
	and pp236(P8[7], X[7], Y[8]);
	and pp237(P8[6], X[6], Y[8]);
	and pp238(P8[5], X[5], Y[8]);
	and pp239(P8[4], X[4], Y[8]);
	and pp240(P8[3], X[3], Y[8]);
	and pp241(P8[2], X[2], Y[8]);
	and pp242(P8[1], X[1], Y[8]);
	and pp243(P8[0], X[0], Y[8]);
	and pp244(sum9[26], X[26], Y[9]);
	and pp245(P9[25], X[25], Y[9]);
	and pp246(P9[24], X[24], Y[9]);
	and pp247(P9[23], X[23], Y[9]);
	and pp248(P9[22], X[22], Y[9]);
	and pp249(P9[21], X[21], Y[9]);
	and pp250(P9[20], X[20], Y[9]);
	and pp251(P9[19], X[19], Y[9]);
	and pp252(P9[18], X[18], Y[9]);
	and pp253(P9[17], X[17], Y[9]);
	and pp254(P9[16], X[16], Y[9]);
	and pp255(P9[15], X[15], Y[9]);
	and pp256(P9[14], X[14], Y[9]);
	and pp257(P9[13], X[13], Y[9]);
	and pp258(P9[12], X[12], Y[9]);
	and pp259(P9[11], X[11], Y[9]);
	and pp260(P9[10], X[10], Y[9]);
	and pp261(P9[9], X[9], Y[9]);
	and pp262(P9[8], X[8], Y[9]);
	and pp263(P9[7], X[7], Y[9]);
	and pp264(P9[6], X[6], Y[9]);
	and pp265(P9[5], X[5], Y[9]);
	and pp266(P9[4], X[4], Y[9]);
	and pp267(P9[3], X[3], Y[9]);
	and pp268(P9[2], X[2], Y[9]);
	and pp269(P9[1], X[1], Y[9]);
	and pp270(P9[0], X[0], Y[9]);
	and pp271(sum10[26], X[26], Y[10]);
	and pp272(P10[25], X[25], Y[10]);
	and pp273(P10[24], X[24], Y[10]);
	and pp274(P10[23], X[23], Y[10]);
	and pp275(P10[22], X[22], Y[10]);
	and pp276(P10[21], X[21], Y[10]);
	and pp277(P10[20], X[20], Y[10]);
	and pp278(P10[19], X[19], Y[10]);
	and pp279(P10[18], X[18], Y[10]);
	and pp280(P10[17], X[17], Y[10]);
	and pp281(P10[16], X[16], Y[10]);
	and pp282(P10[15], X[15], Y[10]);
	and pp283(P10[14], X[14], Y[10]);
	and pp284(P10[13], X[13], Y[10]);
	and pp285(P10[12], X[12], Y[10]);
	and pp286(P10[11], X[11], Y[10]);
	and pp287(P10[10], X[10], Y[10]);
	and pp288(P10[9], X[9], Y[10]);
	and pp289(P10[8], X[8], Y[10]);
	and pp290(P10[7], X[7], Y[10]);
	and pp291(P10[6], X[6], Y[10]);
	and pp292(P10[5], X[5], Y[10]);
	and pp293(P10[4], X[4], Y[10]);
	and pp294(P10[3], X[3], Y[10]);
	and pp295(P10[2], X[2], Y[10]);
	and pp296(P10[1], X[1], Y[10]);
	and pp297(P10[0], X[0], Y[10]);
	and pp298(sum11[26], X[26], Y[11]);
	and pp299(P11[25], X[25], Y[11]);
	and pp300(P11[24], X[24], Y[11]);
	and pp301(P11[23], X[23], Y[11]);
	and pp302(P11[22], X[22], Y[11]);
	and pp303(P11[21], X[21], Y[11]);
	and pp304(P11[20], X[20], Y[11]);
	and pp305(P11[19], X[19], Y[11]);
	and pp306(P11[18], X[18], Y[11]);
	and pp307(P11[17], X[17], Y[11]);
	and pp308(P11[16], X[16], Y[11]);
	and pp309(P11[15], X[15], Y[11]);
	and pp310(P11[14], X[14], Y[11]);
	and pp311(P11[13], X[13], Y[11]);
	and pp312(P11[12], X[12], Y[11]);
	and pp313(P11[11], X[11], Y[11]);
	and pp314(P11[10], X[10], Y[11]);
	and pp315(P11[9], X[9], Y[11]);
	and pp316(P11[8], X[8], Y[11]);
	and pp317(P11[7], X[7], Y[11]);
	and pp318(P11[6], X[6], Y[11]);
	and pp319(P11[5], X[5], Y[11]);
	and pp320(P11[4], X[4], Y[11]);
	and pp321(P11[3], X[3], Y[11]);
	and pp322(P11[2], X[2], Y[11]);
	and pp323(P11[1], X[1], Y[11]);
	and pp324(P11[0], X[0], Y[11]);
	and pp325(sum12[26], X[26], Y[12]);
	and pp326(P12[25], X[25], Y[12]);
	and pp327(P12[24], X[24], Y[12]);
	and pp328(P12[23], X[23], Y[12]);
	and pp329(P12[22], X[22], Y[12]);
	and pp330(P12[21], X[21], Y[12]);
	and pp331(P12[20], X[20], Y[12]);
	and pp332(P12[19], X[19], Y[12]);
	and pp333(P12[18], X[18], Y[12]);
	and pp334(P12[17], X[17], Y[12]);
	and pp335(P12[16], X[16], Y[12]);
	and pp336(P12[15], X[15], Y[12]);
	and pp337(P12[14], X[14], Y[12]);
	and pp338(P12[13], X[13], Y[12]);
	and pp339(P12[12], X[12], Y[12]);
	and pp340(P12[11], X[11], Y[12]);
	and pp341(P12[10], X[10], Y[12]);
	and pp342(P12[9], X[9], Y[12]);
	and pp343(P12[8], X[8], Y[12]);
	and pp344(P12[7], X[7], Y[12]);
	and pp345(P12[6], X[6], Y[12]);
	and pp346(P12[5], X[5], Y[12]);
	and pp347(P12[4], X[4], Y[12]);
	and pp348(P12[3], X[3], Y[12]);
	and pp349(P12[2], X[2], Y[12]);
	and pp350(P12[1], X[1], Y[12]);
	and pp351(P12[0], X[0], Y[12]);
	and pp352(sum13[26], X[26], Y[13]);
	and pp353(P13[25], X[25], Y[13]);
	and pp354(P13[24], X[24], Y[13]);
	and pp355(P13[23], X[23], Y[13]);
	and pp356(P13[22], X[22], Y[13]);
	and pp357(P13[21], X[21], Y[13]);
	and pp358(P13[20], X[20], Y[13]);
	and pp359(P13[19], X[19], Y[13]);
	and pp360(P13[18], X[18], Y[13]);
	and pp361(P13[17], X[17], Y[13]);
	and pp362(P13[16], X[16], Y[13]);
	and pp363(P13[15], X[15], Y[13]);
	and pp364(P13[14], X[14], Y[13]);
	and pp365(P13[13], X[13], Y[13]);
	and pp366(P13[12], X[12], Y[13]);
	and pp367(P13[11], X[11], Y[13]);
	and pp368(P13[10], X[10], Y[13]);
	and pp369(P13[9], X[9], Y[13]);
	and pp370(P13[8], X[8], Y[13]);
	and pp371(P13[7], X[7], Y[13]);
	and pp372(P13[6], X[6], Y[13]);
	and pp373(P13[5], X[5], Y[13]);
	and pp374(P13[4], X[4], Y[13]);
	and pp375(P13[3], X[3], Y[13]);
	and pp376(P13[2], X[2], Y[13]);
	and pp377(P13[1], X[1], Y[13]);
	and pp378(P13[0], X[0], Y[13]);
	and pp379(sum14[26], X[26], Y[14]);
	and pp380(P14[25], X[25], Y[14]);
	and pp381(P14[24], X[24], Y[14]);
	and pp382(P14[23], X[23], Y[14]);
	and pp383(P14[22], X[22], Y[14]);
	and pp384(P14[21], X[21], Y[14]);
	and pp385(P14[20], X[20], Y[14]);
	and pp386(P14[19], X[19], Y[14]);
	and pp387(P14[18], X[18], Y[14]);
	and pp388(P14[17], X[17], Y[14]);
	and pp389(P14[16], X[16], Y[14]);
	and pp390(P14[15], X[15], Y[14]);
	and pp391(P14[14], X[14], Y[14]);
	and pp392(P14[13], X[13], Y[14]);
	and pp393(P14[12], X[12], Y[14]);
	and pp394(P14[11], X[11], Y[14]);
	and pp395(P14[10], X[10], Y[14]);
	and pp396(P14[9], X[9], Y[14]);
	and pp397(P14[8], X[8], Y[14]);
	and pp398(P14[7], X[7], Y[14]);
	and pp399(P14[6], X[6], Y[14]);
	and pp400(P14[5], X[5], Y[14]);
	and pp401(P14[4], X[4], Y[14]);
	and pp402(P14[3], X[3], Y[14]);
	and pp403(P14[2], X[2], Y[14]);
	and pp404(P14[1], X[1], Y[14]);
	and pp405(P14[0], X[0], Y[14]);
	and pp406(sum15[26], X[26], Y[15]);
	and pp407(P15[25], X[25], Y[15]);
	and pp408(P15[24], X[24], Y[15]);
	and pp409(P15[23], X[23], Y[15]);
	and pp410(P15[22], X[22], Y[15]);
	and pp411(P15[21], X[21], Y[15]);
	and pp412(P15[20], X[20], Y[15]);
	and pp413(P15[19], X[19], Y[15]);
	and pp414(P15[18], X[18], Y[15]);
	and pp415(P15[17], X[17], Y[15]);
	and pp416(P15[16], X[16], Y[15]);
	and pp417(P15[15], X[15], Y[15]);
	and pp418(P15[14], X[14], Y[15]);
	and pp419(P15[13], X[13], Y[15]);
	and pp420(P15[12], X[12], Y[15]);
	and pp421(P15[11], X[11], Y[15]);
	and pp422(P15[10], X[10], Y[15]);
	and pp423(P15[9], X[9], Y[15]);
	and pp424(P15[8], X[8], Y[15]);
	and pp425(P15[7], X[7], Y[15]);
	and pp426(P15[6], X[6], Y[15]);
	and pp427(P15[5], X[5], Y[15]);
	and pp428(P15[4], X[4], Y[15]);
	and pp429(P15[3], X[3], Y[15]);
	and pp430(P15[2], X[2], Y[15]);
	and pp431(P15[1], X[1], Y[15]);
	and pp432(P15[0], X[0], Y[15]);
	and pp433(sum16[26], X[26], Y[16]);
	and pp434(P16[25], X[25], Y[16]);
	and pp435(P16[24], X[24], Y[16]);
	and pp436(P16[23], X[23], Y[16]);
	and pp437(P16[22], X[22], Y[16]);
	and pp438(P16[21], X[21], Y[16]);
	and pp439(P16[20], X[20], Y[16]);
	and pp440(P16[19], X[19], Y[16]);
	and pp441(P16[18], X[18], Y[16]);
	and pp442(P16[17], X[17], Y[16]);
	and pp443(P16[16], X[16], Y[16]);
	and pp444(P16[15], X[15], Y[16]);
	and pp445(P16[14], X[14], Y[16]);
	and pp446(P16[13], X[13], Y[16]);
	and pp447(P16[12], X[12], Y[16]);
	and pp448(P16[11], X[11], Y[16]);
	and pp449(P16[10], X[10], Y[16]);
	and pp450(P16[9], X[9], Y[16]);
	and pp451(P16[8], X[8], Y[16]);
	and pp452(P16[7], X[7], Y[16]);
	and pp453(P16[6], X[6], Y[16]);
	and pp454(P16[5], X[5], Y[16]);
	and pp455(P16[4], X[4], Y[16]);
	and pp456(P16[3], X[3], Y[16]);
	and pp457(P16[2], X[2], Y[16]);
	and pp458(P16[1], X[1], Y[16]);
	and pp459(P16[0], X[0], Y[16]);
	and pp460(sum17[26], X[26], Y[17]);
	and pp461(P17[25], X[25], Y[17]);
	and pp462(P17[24], X[24], Y[17]);
	and pp463(P17[23], X[23], Y[17]);
	and pp464(P17[22], X[22], Y[17]);
	and pp465(P17[21], X[21], Y[17]);
	and pp466(P17[20], X[20], Y[17]);
	and pp467(P17[19], X[19], Y[17]);
	and pp468(P17[18], X[18], Y[17]);
	and pp469(P17[17], X[17], Y[17]);
	and pp470(P17[16], X[16], Y[17]);
	and pp471(P17[15], X[15], Y[17]);
	and pp472(P17[14], X[14], Y[17]);
	and pp473(P17[13], X[13], Y[17]);
	and pp474(P17[12], X[12], Y[17]);
	and pp475(P17[11], X[11], Y[17]);
	and pp476(P17[10], X[10], Y[17]);
	and pp477(P17[9], X[9], Y[17]);
	and pp478(P17[8], X[8], Y[17]);
	and pp479(P17[7], X[7], Y[17]);
	and pp480(P17[6], X[6], Y[17]);
	and pp481(P17[5], X[5], Y[17]);
	and pp482(P17[4], X[4], Y[17]);
	and pp483(P17[3], X[3], Y[17]);
	and pp484(P17[2], X[2], Y[17]);
	and pp485(P17[1], X[1], Y[17]);
	and pp486(P17[0], X[0], Y[17]);
	and pp487(sum18[26], X[26], Y[18]);
	and pp488(P18[25], X[25], Y[18]);
	and pp489(P18[24], X[24], Y[18]);
	and pp490(P18[23], X[23], Y[18]);
	and pp491(P18[22], X[22], Y[18]);
	and pp492(P18[21], X[21], Y[18]);
	and pp493(P18[20], X[20], Y[18]);
	and pp494(P18[19], X[19], Y[18]);
	and pp495(P18[18], X[18], Y[18]);
	and pp496(P18[17], X[17], Y[18]);
	and pp497(P18[16], X[16], Y[18]);
	and pp498(P18[15], X[15], Y[18]);
	and pp499(P18[14], X[14], Y[18]);
	and pp500(P18[13], X[13], Y[18]);
	and pp501(P18[12], X[12], Y[18]);
	and pp502(P18[11], X[11], Y[18]);
	and pp503(P18[10], X[10], Y[18]);
	and pp504(P18[9], X[9], Y[18]);
	and pp505(P18[8], X[8], Y[18]);
	and pp506(P18[7], X[7], Y[18]);
	and pp507(P18[6], X[6], Y[18]);
	and pp508(P18[5], X[5], Y[18]);
	and pp509(P18[4], X[4], Y[18]);
	and pp510(P18[3], X[3], Y[18]);
	and pp511(P18[2], X[2], Y[18]);
	and pp512(P18[1], X[1], Y[18]);
	and pp513(P18[0], X[0], Y[18]);
	and pp514(sum19[26], X[26], Y[19]);
	and pp515(P19[25], X[25], Y[19]);
	and pp516(P19[24], X[24], Y[19]);
	and pp517(P19[23], X[23], Y[19]);
	and pp518(P19[22], X[22], Y[19]);
	and pp519(P19[21], X[21], Y[19]);
	and pp520(P19[20], X[20], Y[19]);
	and pp521(P19[19], X[19], Y[19]);
	and pp522(P19[18], X[18], Y[19]);
	and pp523(P19[17], X[17], Y[19]);
	and pp524(P19[16], X[16], Y[19]);
	and pp525(P19[15], X[15], Y[19]);
	and pp526(P19[14], X[14], Y[19]);
	and pp527(P19[13], X[13], Y[19]);
	and pp528(P19[12], X[12], Y[19]);
	and pp529(P19[11], X[11], Y[19]);
	and pp530(P19[10], X[10], Y[19]);
	and pp531(P19[9], X[9], Y[19]);
	and pp532(P19[8], X[8], Y[19]);
	and pp533(P19[7], X[7], Y[19]);
	and pp534(P19[6], X[6], Y[19]);
	and pp535(P19[5], X[5], Y[19]);
	and pp536(P19[4], X[4], Y[19]);
	and pp537(P19[3], X[3], Y[19]);
	and pp538(P19[2], X[2], Y[19]);
	and pp539(P19[1], X[1], Y[19]);
	and pp540(P19[0], X[0], Y[19]);
	and pp541(sum20[26], X[26], Y[20]);
	and pp542(P20[25], X[25], Y[20]);
	and pp543(P20[24], X[24], Y[20]);
	and pp544(P20[23], X[23], Y[20]);
	and pp545(P20[22], X[22], Y[20]);
	and pp546(P20[21], X[21], Y[20]);
	and pp547(P20[20], X[20], Y[20]);
	and pp548(P20[19], X[19], Y[20]);
	and pp549(P20[18], X[18], Y[20]);
	and pp550(P20[17], X[17], Y[20]);
	and pp551(P20[16], X[16], Y[20]);
	and pp552(P20[15], X[15], Y[20]);
	and pp553(P20[14], X[14], Y[20]);
	and pp554(P20[13], X[13], Y[20]);
	and pp555(P20[12], X[12], Y[20]);
	and pp556(P20[11], X[11], Y[20]);
	and pp557(P20[10], X[10], Y[20]);
	and pp558(P20[9], X[9], Y[20]);
	and pp559(P20[8], X[8], Y[20]);
	and pp560(P20[7], X[7], Y[20]);
	and pp561(P20[6], X[6], Y[20]);
	and pp562(P20[5], X[5], Y[20]);
	and pp563(P20[4], X[4], Y[20]);
	and pp564(P20[3], X[3], Y[20]);
	and pp565(P20[2], X[2], Y[20]);
	and pp566(P20[1], X[1], Y[20]);
	and pp567(P20[0], X[0], Y[20]);
	and pp568(sum21[26], X[26], Y[21]);
	and pp569(P21[25], X[25], Y[21]);
	and pp570(P21[24], X[24], Y[21]);
	and pp571(P21[23], X[23], Y[21]);
	and pp572(P21[22], X[22], Y[21]);
	and pp573(P21[21], X[21], Y[21]);
	and pp574(P21[20], X[20], Y[21]);
	and pp575(P21[19], X[19], Y[21]);
	and pp576(P21[18], X[18], Y[21]);
	and pp577(P21[17], X[17], Y[21]);
	and pp578(P21[16], X[16], Y[21]);
	and pp579(P21[15], X[15], Y[21]);
	and pp580(P21[14], X[14], Y[21]);
	and pp581(P21[13], X[13], Y[21]);
	and pp582(P21[12], X[12], Y[21]);
	and pp583(P21[11], X[11], Y[21]);
	and pp584(P21[10], X[10], Y[21]);
	and pp585(P21[9], X[9], Y[21]);
	and pp586(P21[8], X[8], Y[21]);
	and pp587(P21[7], X[7], Y[21]);
	and pp588(P21[6], X[6], Y[21]);
	and pp589(P21[5], X[5], Y[21]);
	and pp590(P21[4], X[4], Y[21]);
	and pp591(P21[3], X[3], Y[21]);
	and pp592(P21[2], X[2], Y[21]);
	and pp593(P21[1], X[1], Y[21]);
	and pp594(P21[0], X[0], Y[21]);
	and pp595(sum22[26], X[26], Y[22]);
	and pp596(P22[25], X[25], Y[22]);
	and pp597(P22[24], X[24], Y[22]);
	and pp598(P22[23], X[23], Y[22]);
	and pp599(P22[22], X[22], Y[22]);
	and pp600(P22[21], X[21], Y[22]);
	and pp601(P22[20], X[20], Y[22]);
	and pp602(P22[19], X[19], Y[22]);
	and pp603(P22[18], X[18], Y[22]);
	and pp604(P22[17], X[17], Y[22]);
	and pp605(P22[16], X[16], Y[22]);
	and pp606(P22[15], X[15], Y[22]);
	and pp607(P22[14], X[14], Y[22]);
	and pp608(P22[13], X[13], Y[22]);
	and pp609(P22[12], X[12], Y[22]);
	and pp610(P22[11], X[11], Y[22]);
	and pp611(P22[10], X[10], Y[22]);
	and pp612(P22[9], X[9], Y[22]);
	and pp613(P22[8], X[8], Y[22]);
	and pp614(P22[7], X[7], Y[22]);
	and pp615(P22[6], X[6], Y[22]);
	and pp616(P22[5], X[5], Y[22]);
	and pp617(P22[4], X[4], Y[22]);
	and pp618(P22[3], X[3], Y[22]);
	and pp619(P22[2], X[2], Y[22]);
	and pp620(P22[1], X[1], Y[22]);
	and pp621(P22[0], X[0], Y[22]);
	and pp622(sum23[26], X[26], Y[23]);
	and pp623(P23[25], X[25], Y[23]);
	and pp624(P23[24], X[24], Y[23]);
	and pp625(P23[23], X[23], Y[23]);
	and pp626(P23[22], X[22], Y[23]);
	and pp627(P23[21], X[21], Y[23]);
	and pp628(P23[20], X[20], Y[23]);
	and pp629(P23[19], X[19], Y[23]);
	and pp630(P23[18], X[18], Y[23]);
	and pp631(P23[17], X[17], Y[23]);
	and pp632(P23[16], X[16], Y[23]);
	and pp633(P23[15], X[15], Y[23]);
	and pp634(P23[14], X[14], Y[23]);
	and pp635(P23[13], X[13], Y[23]);
	and pp636(P23[12], X[12], Y[23]);
	and pp637(P23[11], X[11], Y[23]);
	and pp638(P23[10], X[10], Y[23]);
	and pp639(P23[9], X[9], Y[23]);
	and pp640(P23[8], X[8], Y[23]);
	and pp641(P23[7], X[7], Y[23]);
	and pp642(P23[6], X[6], Y[23]);
	and pp643(P23[5], X[5], Y[23]);
	and pp644(P23[4], X[4], Y[23]);
	and pp645(P23[3], X[3], Y[23]);
	and pp646(P23[2], X[2], Y[23]);
	and pp647(P23[1], X[1], Y[23]);
	and pp648(P23[0], X[0], Y[23]);
	and pp649(sum24[26], X[26], Y[24]);
	and pp650(P24[25], X[25], Y[24]);
	and pp651(P24[24], X[24], Y[24]);
	and pp652(P24[23], X[23], Y[24]);
	and pp653(P24[22], X[22], Y[24]);
	and pp654(P24[21], X[21], Y[24]);
	and pp655(P24[20], X[20], Y[24]);
	and pp656(P24[19], X[19], Y[24]);
	and pp657(P24[18], X[18], Y[24]);
	and pp658(P24[17], X[17], Y[24]);
	and pp659(P24[16], X[16], Y[24]);
	and pp660(P24[15], X[15], Y[24]);
	and pp661(P24[14], X[14], Y[24]);
	and pp662(P24[13], X[13], Y[24]);
	and pp663(P24[12], X[12], Y[24]);
	and pp664(P24[11], X[11], Y[24]);
	and pp665(P24[10], X[10], Y[24]);
	and pp666(P24[9], X[9], Y[24]);
	and pp667(P24[8], X[8], Y[24]);
	and pp668(P24[7], X[7], Y[24]);
	and pp669(P24[6], X[6], Y[24]);
	and pp670(P24[5], X[5], Y[24]);
	and pp671(P24[4], X[4], Y[24]);
	and pp672(P24[3], X[3], Y[24]);
	and pp673(P24[2], X[2], Y[24]);
	and pp674(P24[1], X[1], Y[24]);
	and pp675(P24[0], X[0], Y[24]);
	and pp676(sum25[26], X[26], Y[25]);
	and pp677(P25[25], X[25], Y[25]);
	and pp678(P25[24], X[24], Y[25]);
	and pp679(P25[23], X[23], Y[25]);
	and pp680(P25[22], X[22], Y[25]);
	and pp681(P25[21], X[21], Y[25]);
	and pp682(P25[20], X[20], Y[25]);
	and pp683(P25[19], X[19], Y[25]);
	and pp684(P25[18], X[18], Y[25]);
	and pp685(P25[17], X[17], Y[25]);
	and pp686(P25[16], X[16], Y[25]);
	and pp687(P25[15], X[15], Y[25]);
	and pp688(P25[14], X[14], Y[25]);
	and pp689(P25[13], X[13], Y[25]);
	and pp690(P25[12], X[12], Y[25]);
	and pp691(P25[11], X[11], Y[25]);
	and pp692(P25[10], X[10], Y[25]);
	and pp693(P25[9], X[9], Y[25]);
	and pp694(P25[8], X[8], Y[25]);
	and pp695(P25[7], X[7], Y[25]);
	and pp696(P25[6], X[6], Y[25]);
	and pp697(P25[5], X[5], Y[25]);
	and pp698(P25[4], X[4], Y[25]);
	and pp699(P25[3], X[3], Y[25]);
	and pp700(P25[2], X[2], Y[25]);
	and pp701(P25[1], X[1], Y[25]);
	and pp702(P25[0], X[0], Y[25]);
	and pp703(sum26[26], X[26], Y[26]);
	and pp704(P26[25], X[25], Y[26]);
	and pp705(P26[24], X[24], Y[26]);
	and pp706(P26[23], X[23], Y[26]);
	and pp707(P26[22], X[22], Y[26]);
	and pp708(P26[21], X[21], Y[26]);
	and pp709(P26[20], X[20], Y[26]);
	and pp710(P26[19], X[19], Y[26]);
	and pp711(P26[18], X[18], Y[26]);
	and pp712(P26[17], X[17], Y[26]);
	and pp713(P26[16], X[16], Y[26]);
	and pp714(P26[15], X[15], Y[26]);
	and pp715(P26[14], X[14], Y[26]);
	and pp716(P26[13], X[13], Y[26]);
	and pp717(P26[12], X[12], Y[26]);
	and pp718(P26[11], X[11], Y[26]);
	and pp719(P26[10], X[10], Y[26]);
	and pp720(P26[9], X[9], Y[26]);
	and pp721(P26[8], X[8], Y[26]);
	and pp722(P26[7], X[7], Y[26]);
	and pp723(P26[6], X[6], Y[26]);
	and pp724(P26[5], X[5], Y[26]);
	and pp725(P26[4], X[4], Y[26]);
	and pp726(P26[3], X[3], Y[26]);
	and pp727(P26[2], X[2], Y[26]);
	and pp728(P26[1], X[1], Y[26]);
	and pp729(P26[0], X[0], Y[26]);

	// Array Reduction
	half_adder  HA1(carry1[25],sum1[25],P1[25],P0[26]);
	half_adder  HA2(carry1[24],sum1[24],P1[24],P0[25]);
	half_adder  HA3(carry1[23],sum1[23],P1[23],P0[24]);
	half_adder  HA4(carry1[22],sum1[22],P1[22],P0[23]);
	half_adder  HA5(carry1[21],sum1[21],P1[21],P0[22]);
	half_adder  HA6(carry1[20],sum1[20],P1[20],P0[21]);
	half_adder  HA7(carry1[19],sum1[19],P1[19],P0[20]);
	half_adder  HA8(carry1[18],sum1[18],P1[18],P0[19]);
	half_adder  HA9(carry1[17],sum1[17],P1[17],P0[18]);
	half_adder  HA10(carry1[16],sum1[16],P1[16],P0[17]);
	half_adder  HA11(carry1[15],sum1[15],P1[15],P0[16]);
	half_adder  HA12(carry1[14],sum1[14],P1[14],P0[15]);
	half_adder  HA13(carry1[13],sum1[13],P1[13],P0[14]);
	half_adder  HA14(carry1[12],sum1[12],P1[12],P0[13]);
	half_adder  HA15(carry1[11],sum1[11],P1[11],P0[12]);
	half_adder  HA16(carry1[10],sum1[10],P1[10],P0[11]);
	half_adder  HA17(carry1[9],sum1[9],P1[9],P0[10]);
	half_adder  HA18(carry1[8],sum1[8],P1[8],P0[9]);
	half_adder  HA19(carry1[7],sum1[7],P1[7],P0[8]);
	half_adder  HA20(carry1[6],sum1[6],P1[6],P0[7]);
	half_adder  HA21(carry1[5],sum1[5],P1[5],P0[6]);
	half_adder  HA22(carry1[4],sum1[4],P1[4],P0[5]);
	half_adder  HA23(carry1[3],sum1[3],P1[3],P0[4]);
	half_adder  HA24(carry1[2],sum1[2],P1[2],P0[3]);
	half_adder  HA25(carry1[1],sum1[1],P1[1],P0[2]);
	half_adder  HA26(carry1[0],sum1[0],P1[0],P0[1]);
	full_adder  FA1(carry2[25],sum2[25],P2[25],sum1[26],carry1[25]);
	full_adder  FA2(carry2[24],sum2[24],P2[24],sum1[25],carry1[24]);
	full_adder  FA3(carry2[23],sum2[23],P2[23],sum1[24],carry1[23]);
	full_adder  FA4(carry2[22],sum2[22],P2[22],sum1[23],carry1[22]);
	full_adder  FA5(carry2[21],sum2[21],P2[21],sum1[22],carry1[21]);
	full_adder  FA6(carry2[20],sum2[20],P2[20],sum1[21],carry1[20]);
	full_adder  FA7(carry2[19],sum2[19],P2[19],sum1[20],carry1[19]);
	full_adder  FA8(carry2[18],sum2[18],P2[18],sum1[19],carry1[18]);
	full_adder  FA9(carry2[17],sum2[17],P2[17],sum1[18],carry1[17]);
	full_adder  FA10(carry2[16],sum2[16],P2[16],sum1[17],carry1[16]);
	full_adder  FA11(carry2[15],sum2[15],P2[15],sum1[16],carry1[15]);
	full_adder  FA12(carry2[14],sum2[14],P2[14],sum1[15],carry1[14]);
	full_adder  FA13(carry2[13],sum2[13],P2[13],sum1[14],carry1[13]);
	full_adder  FA14(carry2[12],sum2[12],P2[12],sum1[13],carry1[12]);
	full_adder  FA15(carry2[11],sum2[11],P2[11],sum1[12],carry1[11]);
	full_adder  FA16(carry2[10],sum2[10],P2[10],sum1[11],carry1[10]);
	full_adder  FA17(carry2[9],sum2[9],P2[9],sum1[10],carry1[9]);
	full_adder  FA18(carry2[8],sum2[8],P2[8],sum1[9],carry1[8]);
	full_adder  FA19(carry2[7],sum2[7],P2[7],sum1[8],carry1[7]);
	full_adder  FA20(carry2[6],sum2[6],P2[6],sum1[7],carry1[6]);
	full_adder  FA21(carry2[5],sum2[5],P2[5],sum1[6],carry1[5]);
	full_adder  FA22(carry2[4],sum2[4],P2[4],sum1[5],carry1[4]);
	full_adder  FA23(carry2[3],sum2[3],P2[3],sum1[4],carry1[3]);
	full_adder  FA24(carry2[2],sum2[2],P2[2],sum1[3],carry1[2]);
	full_adder  FA25(carry2[1],sum2[1],P2[1],sum1[2],carry1[1]);
	full_adder  FA26(carry2[0],sum2[0],P2[0],sum1[1],carry1[0]);
	full_adder  FA27(carry3[25],sum3[25],P3[25],sum2[26],carry2[25]);
	full_adder  FA28(carry3[24],sum3[24],P3[24],sum2[25],carry2[24]);
	full_adder  FA29(carry3[23],sum3[23],P3[23],sum2[24],carry2[23]);
	full_adder  FA30(carry3[22],sum3[22],P3[22],sum2[23],carry2[22]);
	full_adder  FA31(carry3[21],sum3[21],P3[21],sum2[22],carry2[21]);
	full_adder  FA32(carry3[20],sum3[20],P3[20],sum2[21],carry2[20]);
	full_adder  FA33(carry3[19],sum3[19],P3[19],sum2[20],carry2[19]);
	full_adder  FA34(carry3[18],sum3[18],P3[18],sum2[19],carry2[18]);
	full_adder  FA35(carry3[17],sum3[17],P3[17],sum2[18],carry2[17]);
	full_adder  FA36(carry3[16],sum3[16],P3[16],sum2[17],carry2[16]);
	full_adder  FA37(carry3[15],sum3[15],P3[15],sum2[16],carry2[15]);
	full_adder  FA38(carry3[14],sum3[14],P3[14],sum2[15],carry2[14]);
	full_adder  FA39(carry3[13],sum3[13],P3[13],sum2[14],carry2[13]);
	full_adder  FA40(carry3[12],sum3[12],P3[12],sum2[13],carry2[12]);
	full_adder  FA41(carry3[11],sum3[11],P3[11],sum2[12],carry2[11]);
	full_adder  FA42(carry3[10],sum3[10],P3[10],sum2[11],carry2[10]);
	full_adder  FA43(carry3[9],sum3[9],P3[9],sum2[10],carry2[9]);
	full_adder  FA44(carry3[8],sum3[8],P3[8],sum2[9],carry2[8]);
	full_adder  FA45(carry3[7],sum3[7],P3[7],sum2[8],carry2[7]);
	full_adder  FA46(carry3[6],sum3[6],P3[6],sum2[7],carry2[6]);
	full_adder  FA47(carry3[5],sum3[5],P3[5],sum2[6],carry2[5]);
	full_adder  FA48(carry3[4],sum3[4],P3[4],sum2[5],carry2[4]);
	full_adder  FA49(carry3[3],sum3[3],P3[3],sum2[4],carry2[3]);
	full_adder  FA50(carry3[2],sum3[2],P3[2],sum2[3],carry2[2]);
	full_adder  FA51(carry3[1],sum3[1],P3[1],sum2[2],carry2[1]);
	full_adder  FA52(carry3[0],sum3[0],P3[0],sum2[1],carry2[0]);
	full_adder  FA53(carry4[25],sum4[25],P4[25],sum3[26],carry3[25]);
	full_adder  FA54(carry4[24],sum4[24],P4[24],sum3[25],carry3[24]);
	full_adder  FA55(carry4[23],sum4[23],P4[23],sum3[24],carry3[23]);
	full_adder  FA56(carry4[22],sum4[22],P4[22],sum3[23],carry3[22]);
	full_adder  FA57(carry4[21],sum4[21],P4[21],sum3[22],carry3[21]);
	full_adder  FA58(carry4[20],sum4[20],P4[20],sum3[21],carry3[20]);
	full_adder  FA59(carry4[19],sum4[19],P4[19],sum3[20],carry3[19]);
	full_adder  FA60(carry4[18],sum4[18],P4[18],sum3[19],carry3[18]);
	full_adder  FA61(carry4[17],sum4[17],P4[17],sum3[18],carry3[17]);
	full_adder  FA62(carry4[16],sum4[16],P4[16],sum3[17],carry3[16]);
	full_adder  FA63(carry4[15],sum4[15],P4[15],sum3[16],carry3[15]);
	full_adder  FA64(carry4[14],sum4[14],P4[14],sum3[15],carry3[14]);
	full_adder  FA65(carry4[13],sum4[13],P4[13],sum3[14],carry3[13]);
	full_adder  FA66(carry4[12],sum4[12],P4[12],sum3[13],carry3[12]);
	full_adder  FA67(carry4[11],sum4[11],P4[11],sum3[12],carry3[11]);
	full_adder  FA68(carry4[10],sum4[10],P4[10],sum3[11],carry3[10]);
	full_adder  FA69(carry4[9],sum4[9],P4[9],sum3[10],carry3[9]);
	full_adder  FA70(carry4[8],sum4[8],P4[8],sum3[9],carry3[8]);
	full_adder  FA71(carry4[7],sum4[7],P4[7],sum3[8],carry3[7]);
	full_adder  FA72(carry4[6],sum4[6],P4[6],sum3[7],carry3[6]);
	full_adder  FA73(carry4[5],sum4[5],P4[5],sum3[6],carry3[5]);
	full_adder  FA74(carry4[4],sum4[4],P4[4],sum3[5],carry3[4]);
	full_adder  FA75(carry4[3],sum4[3],P4[3],sum3[4],carry3[3]);
	full_adder  FA76(carry4[2],sum4[2],P4[2],sum3[3],carry3[2]);
	full_adder  FA77(carry4[1],sum4[1],P4[1],sum3[2],carry3[1]);
	full_adder  FA78(carry4[0],sum4[0],P4[0],sum3[1],carry3[0]);
	full_adder  FA79(carry5[25],sum5[25],P5[25],sum4[26],carry4[25]);
	full_adder  FA80(carry5[24],sum5[24],P5[24],sum4[25],carry4[24]);
	full_adder  FA81(carry5[23],sum5[23],P5[23],sum4[24],carry4[23]);
	full_adder  FA82(carry5[22],sum5[22],P5[22],sum4[23],carry4[22]);
	full_adder  FA83(carry5[21],sum5[21],P5[21],sum4[22],carry4[21]);
	full_adder  FA84(carry5[20],sum5[20],P5[20],sum4[21],carry4[20]);
	full_adder  FA85(carry5[19],sum5[19],P5[19],sum4[20],carry4[19]);
	full_adder  FA86(carry5[18],sum5[18],P5[18],sum4[19],carry4[18]);
	full_adder  FA87(carry5[17],sum5[17],P5[17],sum4[18],carry4[17]);
	full_adder  FA88(carry5[16],sum5[16],P5[16],sum4[17],carry4[16]);
	full_adder  FA89(carry5[15],sum5[15],P5[15],sum4[16],carry4[15]);
	full_adder  FA90(carry5[14],sum5[14],P5[14],sum4[15],carry4[14]);
	full_adder  FA91(carry5[13],sum5[13],P5[13],sum4[14],carry4[13]);
	full_adder  FA92(carry5[12],sum5[12],P5[12],sum4[13],carry4[12]);
	full_adder  FA93(carry5[11],sum5[11],P5[11],sum4[12],carry4[11]);
	full_adder  FA94(carry5[10],sum5[10],P5[10],sum4[11],carry4[10]);
	full_adder  FA95(carry5[9],sum5[9],P5[9],sum4[10],carry4[9]);
	full_adder  FA96(carry5[8],sum5[8],P5[8],sum4[9],carry4[8]);
	full_adder  FA97(carry5[7],sum5[7],P5[7],sum4[8],carry4[7]);
	full_adder  FA98(carry5[6],sum5[6],P5[6],sum4[7],carry4[6]);
	full_adder  FA99(carry5[5],sum5[5],P5[5],sum4[6],carry4[5]);
	full_adder  FA100(carry5[4],sum5[4],P5[4],sum4[5],carry4[4]);
	full_adder  FA101(carry5[3],sum5[3],P5[3],sum4[4],carry4[3]);
	full_adder  FA102(carry5[2],sum5[2],P5[2],sum4[3],carry4[2]);
	full_adder  FA103(carry5[1],sum5[1],P5[1],sum4[2],carry4[1]);
	full_adder  FA104(carry5[0],sum5[0],P5[0],sum4[1],carry4[0]);
	full_adder  FA105(carry6[25],sum6[25],P6[25],sum5[26],carry5[25]);
	full_adder  FA106(carry6[24],sum6[24],P6[24],sum5[25],carry5[24]);
	full_adder  FA107(carry6[23],sum6[23],P6[23],sum5[24],carry5[23]);
	full_adder  FA108(carry6[22],sum6[22],P6[22],sum5[23],carry5[22]);
	full_adder  FA109(carry6[21],sum6[21],P6[21],sum5[22],carry5[21]);
	full_adder  FA110(carry6[20],sum6[20],P6[20],sum5[21],carry5[20]);
	full_adder  FA111(carry6[19],sum6[19],P6[19],sum5[20],carry5[19]);
	full_adder  FA112(carry6[18],sum6[18],P6[18],sum5[19],carry5[18]);
	full_adder  FA113(carry6[17],sum6[17],P6[17],sum5[18],carry5[17]);
	full_adder  FA114(carry6[16],sum6[16],P6[16],sum5[17],carry5[16]);
	full_adder  FA115(carry6[15],sum6[15],P6[15],sum5[16],carry5[15]);
	full_adder  FA116(carry6[14],sum6[14],P6[14],sum5[15],carry5[14]);
	full_adder  FA117(carry6[13],sum6[13],P6[13],sum5[14],carry5[13]);
	full_adder  FA118(carry6[12],sum6[12],P6[12],sum5[13],carry5[12]);
	full_adder  FA119(carry6[11],sum6[11],P6[11],sum5[12],carry5[11]);
	full_adder  FA120(carry6[10],sum6[10],P6[10],sum5[11],carry5[10]);
	full_adder  FA121(carry6[9],sum6[9],P6[9],sum5[10],carry5[9]);
	full_adder  FA122(carry6[8],sum6[8],P6[8],sum5[9],carry5[8]);
	full_adder  FA123(carry6[7],sum6[7],P6[7],sum5[8],carry5[7]);
	full_adder  FA124(carry6[6],sum6[6],P6[6],sum5[7],carry5[6]);
	full_adder  FA125(carry6[5],sum6[5],P6[5],sum5[6],carry5[5]);
	full_adder  FA126(carry6[4],sum6[4],P6[4],sum5[5],carry5[4]);
	full_adder  FA127(carry6[3],sum6[3],P6[3],sum5[4],carry5[3]);
	full_adder  FA128(carry6[2],sum6[2],P6[2],sum5[3],carry5[2]);
	full_adder  FA129(carry6[1],sum6[1],P6[1],sum5[2],carry5[1]);
	full_adder  FA130(carry6[0],sum6[0],P6[0],sum5[1],carry5[0]);
	full_adder  FA131(carry7[25],sum7[25],P7[25],sum6[26],carry6[25]);
	full_adder  FA132(carry7[24],sum7[24],P7[24],sum6[25],carry6[24]);
	full_adder  FA133(carry7[23],sum7[23],P7[23],sum6[24],carry6[23]);
	full_adder  FA134(carry7[22],sum7[22],P7[22],sum6[23],carry6[22]);
	full_adder  FA135(carry7[21],sum7[21],P7[21],sum6[22],carry6[21]);
	full_adder  FA136(carry7[20],sum7[20],P7[20],sum6[21],carry6[20]);
	full_adder  FA137(carry7[19],sum7[19],P7[19],sum6[20],carry6[19]);
	full_adder  FA138(carry7[18],sum7[18],P7[18],sum6[19],carry6[18]);
	full_adder  FA139(carry7[17],sum7[17],P7[17],sum6[18],carry6[17]);
	full_adder  FA140(carry7[16],sum7[16],P7[16],sum6[17],carry6[16]);
	full_adder  FA141(carry7[15],sum7[15],P7[15],sum6[16],carry6[15]);
	full_adder  FA142(carry7[14],sum7[14],P7[14],sum6[15],carry6[14]);
	full_adder  FA143(carry7[13],sum7[13],P7[13],sum6[14],carry6[13]);
	full_adder  FA144(carry7[12],sum7[12],P7[12],sum6[13],carry6[12]);
	full_adder  FA145(carry7[11],sum7[11],P7[11],sum6[12],carry6[11]);
	full_adder  FA146(carry7[10],sum7[10],P7[10],sum6[11],carry6[10]);
	full_adder  FA147(carry7[9],sum7[9],P7[9],sum6[10],carry6[9]);
	full_adder  FA148(carry7[8],sum7[8],P7[8],sum6[9],carry6[8]);
	full_adder  FA149(carry7[7],sum7[7],P7[7],sum6[8],carry6[7]);
	full_adder  FA150(carry7[6],sum7[6],P7[6],sum6[7],carry6[6]);
	full_adder  FA151(carry7[5],sum7[5],P7[5],sum6[6],carry6[5]);
	full_adder  FA152(carry7[4],sum7[4],P7[4],sum6[5],carry6[4]);
	full_adder  FA153(carry7[3],sum7[3],P7[3],sum6[4],carry6[3]);
	full_adder  FA154(carry7[2],sum7[2],P7[2],sum6[3],carry6[2]);
	full_adder  FA155(carry7[1],sum7[1],P7[1],sum6[2],carry6[1]);
	full_adder  FA156(carry7[0],sum7[0],P7[0],sum6[1],carry6[0]);
	full_adder  FA157(carry8[25],sum8[25],P8[25],sum7[26],carry7[25]);
	full_adder  FA158(carry8[24],sum8[24],P8[24],sum7[25],carry7[24]);
	full_adder  FA159(carry8[23],sum8[23],P8[23],sum7[24],carry7[23]);
	full_adder  FA160(carry8[22],sum8[22],P8[22],sum7[23],carry7[22]);
	full_adder  FA161(carry8[21],sum8[21],P8[21],sum7[22],carry7[21]);
	full_adder  FA162(carry8[20],sum8[20],P8[20],sum7[21],carry7[20]);
	full_adder  FA163(carry8[19],sum8[19],P8[19],sum7[20],carry7[19]);
	full_adder  FA164(carry8[18],sum8[18],P8[18],sum7[19],carry7[18]);
	full_adder  FA165(carry8[17],sum8[17],P8[17],sum7[18],carry7[17]);
	full_adder  FA166(carry8[16],sum8[16],P8[16],sum7[17],carry7[16]);
	full_adder  FA167(carry8[15],sum8[15],P8[15],sum7[16],carry7[15]);
	full_adder  FA168(carry8[14],sum8[14],P8[14],sum7[15],carry7[14]);
	full_adder  FA169(carry8[13],sum8[13],P8[13],sum7[14],carry7[13]);
	full_adder  FA170(carry8[12],sum8[12],P8[12],sum7[13],carry7[12]);
	full_adder  FA171(carry8[11],sum8[11],P8[11],sum7[12],carry7[11]);
	full_adder  FA172(carry8[10],sum8[10],P8[10],sum7[11],carry7[10]);
	full_adder  FA173(carry8[9],sum8[9],P8[9],sum7[10],carry7[9]);
	full_adder  FA174(carry8[8],sum8[8],P8[8],sum7[9],carry7[8]);
	full_adder  FA175(carry8[7],sum8[7],P8[7],sum7[8],carry7[7]);
	full_adder  FA176(carry8[6],sum8[6],P8[6],sum7[7],carry7[6]);
	full_adder  FA177(carry8[5],sum8[5],P8[5],sum7[6],carry7[5]);
	full_adder  FA178(carry8[4],sum8[4],P8[4],sum7[5],carry7[4]);
	full_adder  FA179(carry8[3],sum8[3],P8[3],sum7[4],carry7[3]);
	full_adder  FA180(carry8[2],sum8[2],P8[2],sum7[3],carry7[2]);
	full_adder  FA181(carry8[1],sum8[1],P8[1],sum7[2],carry7[1]);
	full_adder  FA182(carry8[0],sum8[0],P8[0],sum7[1],carry7[0]);
	full_adder  FA183(carry9[25],sum9[25],P9[25],sum8[26],carry8[25]);
	full_adder  FA184(carry9[24],sum9[24],P9[24],sum8[25],carry8[24]);
	full_adder  FA185(carry9[23],sum9[23],P9[23],sum8[24],carry8[23]);
	full_adder  FA186(carry9[22],sum9[22],P9[22],sum8[23],carry8[22]);
	full_adder  FA187(carry9[21],sum9[21],P9[21],sum8[22],carry8[21]);
	full_adder  FA188(carry9[20],sum9[20],P9[20],sum8[21],carry8[20]);
	full_adder  FA189(carry9[19],sum9[19],P9[19],sum8[20],carry8[19]);
	full_adder  FA190(carry9[18],sum9[18],P9[18],sum8[19],carry8[18]);
	full_adder  FA191(carry9[17],sum9[17],P9[17],sum8[18],carry8[17]);
	full_adder  FA192(carry9[16],sum9[16],P9[16],sum8[17],carry8[16]);
	full_adder  FA193(carry9[15],sum9[15],P9[15],sum8[16],carry8[15]);
	full_adder  FA194(carry9[14],sum9[14],P9[14],sum8[15],carry8[14]);
	full_adder  FA195(carry9[13],sum9[13],P9[13],sum8[14],carry8[13]);
	full_adder  FA196(carry9[12],sum9[12],P9[12],sum8[13],carry8[12]);
	full_adder  FA197(carry9[11],sum9[11],P9[11],sum8[12],carry8[11]);
	full_adder  FA198(carry9[10],sum9[10],P9[10],sum8[11],carry8[10]);
	full_adder  FA199(carry9[9],sum9[9],P9[9],sum8[10],carry8[9]);
	full_adder  FA200(carry9[8],sum9[8],P9[8],sum8[9],carry8[8]);
	full_adder  FA201(carry9[7],sum9[7],P9[7],sum8[8],carry8[7]);
	full_adder  FA202(carry9[6],sum9[6],P9[6],sum8[7],carry8[6]);
	full_adder  FA203(carry9[5],sum9[5],P9[5],sum8[6],carry8[5]);
	full_adder  FA204(carry9[4],sum9[4],P9[4],sum8[5],carry8[4]);
	full_adder  FA205(carry9[3],sum9[3],P9[3],sum8[4],carry8[3]);
	full_adder  FA206(carry9[2],sum9[2],P9[2],sum8[3],carry8[2]);
	full_adder  FA207(carry9[1],sum9[1],P9[1],sum8[2],carry8[1]);
	full_adder  FA208(carry9[0],sum9[0],P9[0],sum8[1],carry8[0]);
	full_adder  FA209(carry10[25],sum10[25],P10[25],sum9[26],carry9[25]);
	full_adder  FA210(carry10[24],sum10[24],P10[24],sum9[25],carry9[24]);
	full_adder  FA211(carry10[23],sum10[23],P10[23],sum9[24],carry9[23]);
	full_adder  FA212(carry10[22],sum10[22],P10[22],sum9[23],carry9[22]);
	full_adder  FA213(carry10[21],sum10[21],P10[21],sum9[22],carry9[21]);
	full_adder  FA214(carry10[20],sum10[20],P10[20],sum9[21],carry9[20]);
	full_adder  FA215(carry10[19],sum10[19],P10[19],sum9[20],carry9[19]);
	full_adder  FA216(carry10[18],sum10[18],P10[18],sum9[19],carry9[18]);
	full_adder  FA217(carry10[17],sum10[17],P10[17],sum9[18],carry9[17]);
	full_adder  FA218(carry10[16],sum10[16],P10[16],sum9[17],carry9[16]);
	full_adder  FA219(carry10[15],sum10[15],P10[15],sum9[16],carry9[15]);
	full_adder  FA220(carry10[14],sum10[14],P10[14],sum9[15],carry9[14]);
	full_adder  FA221(carry10[13],sum10[13],P10[13],sum9[14],carry9[13]);
	full_adder  FA222(carry10[12],sum10[12],P10[12],sum9[13],carry9[12]);
	full_adder  FA223(carry10[11],sum10[11],P10[11],sum9[12],carry9[11]);
	full_adder  FA224(carry10[10],sum10[10],P10[10],sum9[11],carry9[10]);
	full_adder  FA225(carry10[9],sum10[9],P10[9],sum9[10],carry9[9]);
	full_adder  FA226(carry10[8],sum10[8],P10[8],sum9[9],carry9[8]);
	full_adder  FA227(carry10[7],sum10[7],P10[7],sum9[8],carry9[7]);
	full_adder  FA228(carry10[6],sum10[6],P10[6],sum9[7],carry9[6]);
	full_adder  FA229(carry10[5],sum10[5],P10[5],sum9[6],carry9[5]);
	full_adder  FA230(carry10[4],sum10[4],P10[4],sum9[5],carry9[4]);
	full_adder  FA231(carry10[3],sum10[3],P10[3],sum9[4],carry9[3]);
	full_adder  FA232(carry10[2],sum10[2],P10[2],sum9[3],carry9[2]);
	full_adder  FA233(carry10[1],sum10[1],P10[1],sum9[2],carry9[1]);
	full_adder  FA234(carry10[0],sum10[0],P10[0],sum9[1],carry9[0]);
	full_adder  FA235(carry11[25],sum11[25],P11[25],sum10[26],carry10[25]);
	full_adder  FA236(carry11[24],sum11[24],P11[24],sum10[25],carry10[24]);
	full_adder  FA237(carry11[23],sum11[23],P11[23],sum10[24],carry10[23]);
	full_adder  FA238(carry11[22],sum11[22],P11[22],sum10[23],carry10[22]);
	full_adder  FA239(carry11[21],sum11[21],P11[21],sum10[22],carry10[21]);
	full_adder  FA240(carry11[20],sum11[20],P11[20],sum10[21],carry10[20]);
	full_adder  FA241(carry11[19],sum11[19],P11[19],sum10[20],carry10[19]);
	full_adder  FA242(carry11[18],sum11[18],P11[18],sum10[19],carry10[18]);
	full_adder  FA243(carry11[17],sum11[17],P11[17],sum10[18],carry10[17]);
	full_adder  FA244(carry11[16],sum11[16],P11[16],sum10[17],carry10[16]);
	full_adder  FA245(carry11[15],sum11[15],P11[15],sum10[16],carry10[15]);
	full_adder  FA246(carry11[14],sum11[14],P11[14],sum10[15],carry10[14]);
	full_adder  FA247(carry11[13],sum11[13],P11[13],sum10[14],carry10[13]);
	full_adder  FA248(carry11[12],sum11[12],P11[12],sum10[13],carry10[12]);
	full_adder  FA249(carry11[11],sum11[11],P11[11],sum10[12],carry10[11]);
	full_adder  FA250(carry11[10],sum11[10],P11[10],sum10[11],carry10[10]);
	full_adder  FA251(carry11[9],sum11[9],P11[9],sum10[10],carry10[9]);
	full_adder  FA252(carry11[8],sum11[8],P11[8],sum10[9],carry10[8]);
	full_adder  FA253(carry11[7],sum11[7],P11[7],sum10[8],carry10[7]);
	full_adder  FA254(carry11[6],sum11[6],P11[6],sum10[7],carry10[6]);
	full_adder  FA255(carry11[5],sum11[5],P11[5],sum10[6],carry10[5]);
	full_adder  FA256(carry11[4],sum11[4],P11[4],sum10[5],carry10[4]);
	full_adder  FA257(carry11[3],sum11[3],P11[3],sum10[4],carry10[3]);
	full_adder  FA258(carry11[2],sum11[2],P11[2],sum10[3],carry10[2]);
	full_adder  FA259(carry11[1],sum11[1],P11[1],sum10[2],carry10[1]);
	full_adder  FA260(carry11[0],sum11[0],P11[0],sum10[1],carry10[0]);
	full_adder  FA261(carry12[25],sum12[25],P12[25],sum11[26],carry11[25]);
	full_adder  FA262(carry12[24],sum12[24],P12[24],sum11[25],carry11[24]);
	full_adder  FA263(carry12[23],sum12[23],P12[23],sum11[24],carry11[23]);
	full_adder  FA264(carry12[22],sum12[22],P12[22],sum11[23],carry11[22]);
	full_adder  FA265(carry12[21],sum12[21],P12[21],sum11[22],carry11[21]);
	full_adder  FA266(carry12[20],sum12[20],P12[20],sum11[21],carry11[20]);
	full_adder  FA267(carry12[19],sum12[19],P12[19],sum11[20],carry11[19]);
	full_adder  FA268(carry12[18],sum12[18],P12[18],sum11[19],carry11[18]);
	full_adder  FA269(carry12[17],sum12[17],P12[17],sum11[18],carry11[17]);
	full_adder  FA270(carry12[16],sum12[16],P12[16],sum11[17],carry11[16]);
	full_adder  FA271(carry12[15],sum12[15],P12[15],sum11[16],carry11[15]);
	full_adder  FA272(carry12[14],sum12[14],P12[14],sum11[15],carry11[14]);
	full_adder  FA273(carry12[13],sum12[13],P12[13],sum11[14],carry11[13]);
	full_adder  FA274(carry12[12],sum12[12],P12[12],sum11[13],carry11[12]);
	full_adder  FA275(carry12[11],sum12[11],P12[11],sum11[12],carry11[11]);
	full_adder  FA276(carry12[10],sum12[10],P12[10],sum11[11],carry11[10]);
	full_adder  FA277(carry12[9],sum12[9],P12[9],sum11[10],carry11[9]);
	full_adder  FA278(carry12[8],sum12[8],P12[8],sum11[9],carry11[8]);
	full_adder  FA279(carry12[7],sum12[7],P12[7],sum11[8],carry11[7]);
	full_adder  FA280(carry12[6],sum12[6],P12[6],sum11[7],carry11[6]);
	full_adder  FA281(carry12[5],sum12[5],P12[5],sum11[6],carry11[5]);
	full_adder  FA282(carry12[4],sum12[4],P12[4],sum11[5],carry11[4]);
	full_adder  FA283(carry12[3],sum12[3],P12[3],sum11[4],carry11[3]);
	full_adder  FA284(carry12[2],sum12[2],P12[2],sum11[3],carry11[2]);
	full_adder  FA285(carry12[1],sum12[1],P12[1],sum11[2],carry11[1]);
	full_adder  FA286(carry12[0],sum12[0],P12[0],sum11[1],carry11[0]);
	full_adder  FA287(carry13[25],sum13[25],P13[25],sum12[26],carry12[25]);
	full_adder  FA288(carry13[24],sum13[24],P13[24],sum12[25],carry12[24]);
	full_adder  FA289(carry13[23],sum13[23],P13[23],sum12[24],carry12[23]);
	full_adder  FA290(carry13[22],sum13[22],P13[22],sum12[23],carry12[22]);
	full_adder  FA291(carry13[21],sum13[21],P13[21],sum12[22],carry12[21]);
	full_adder  FA292(carry13[20],sum13[20],P13[20],sum12[21],carry12[20]);
	full_adder  FA293(carry13[19],sum13[19],P13[19],sum12[20],carry12[19]);
	full_adder  FA294(carry13[18],sum13[18],P13[18],sum12[19],carry12[18]);
	full_adder  FA295(carry13[17],sum13[17],P13[17],sum12[18],carry12[17]);
	full_adder  FA296(carry13[16],sum13[16],P13[16],sum12[17],carry12[16]);
	full_adder  FA297(carry13[15],sum13[15],P13[15],sum12[16],carry12[15]);
	full_adder  FA298(carry13[14],sum13[14],P13[14],sum12[15],carry12[14]);
	full_adder  FA299(carry13[13],sum13[13],P13[13],sum12[14],carry12[13]);
	full_adder  FA300(carry13[12],sum13[12],P13[12],sum12[13],carry12[12]);
	full_adder  FA301(carry13[11],sum13[11],P13[11],sum12[12],carry12[11]);
	full_adder  FA302(carry13[10],sum13[10],P13[10],sum12[11],carry12[10]);
	full_adder  FA303(carry13[9],sum13[9],P13[9],sum12[10],carry12[9]);
	full_adder  FA304(carry13[8],sum13[8],P13[8],sum12[9],carry12[8]);
	full_adder  FA305(carry13[7],sum13[7],P13[7],sum12[8],carry12[7]);
	full_adder  FA306(carry13[6],sum13[6],P13[6],sum12[7],carry12[6]);
	full_adder  FA307(carry13[5],sum13[5],P13[5],sum12[6],carry12[5]);
	full_adder  FA308(carry13[4],sum13[4],P13[4],sum12[5],carry12[4]);
	full_adder  FA309(carry13[3],sum13[3],P13[3],sum12[4],carry12[3]);
	full_adder  FA310(carry13[2],sum13[2],P13[2],sum12[3],carry12[2]);
	full_adder  FA311(carry13[1],sum13[1],P13[1],sum12[2],carry12[1]);
	full_adder  FA312(carry13[0],sum13[0],P13[0],sum12[1],carry12[0]);
	full_adder  FA313(carry14[25],sum14[25],P14[25],sum13[26],carry13[25]);
	full_adder  FA314(carry14[24],sum14[24],P14[24],sum13[25],carry13[24]);
	full_adder  FA315(carry14[23],sum14[23],P14[23],sum13[24],carry13[23]);
	full_adder  FA316(carry14[22],sum14[22],P14[22],sum13[23],carry13[22]);
	full_adder  FA317(carry14[21],sum14[21],P14[21],sum13[22],carry13[21]);
	full_adder  FA318(carry14[20],sum14[20],P14[20],sum13[21],carry13[20]);
	full_adder  FA319(carry14[19],sum14[19],P14[19],sum13[20],carry13[19]);
	full_adder  FA320(carry14[18],sum14[18],P14[18],sum13[19],carry13[18]);
	full_adder  FA321(carry14[17],sum14[17],P14[17],sum13[18],carry13[17]);
	full_adder  FA322(carry14[16],sum14[16],P14[16],sum13[17],carry13[16]);
	full_adder  FA323(carry14[15],sum14[15],P14[15],sum13[16],carry13[15]);
	full_adder  FA324(carry14[14],sum14[14],P14[14],sum13[15],carry13[14]);
	full_adder  FA325(carry14[13],sum14[13],P14[13],sum13[14],carry13[13]);
	full_adder  FA326(carry14[12],sum14[12],P14[12],sum13[13],carry13[12]);
	full_adder  FA327(carry14[11],sum14[11],P14[11],sum13[12],carry13[11]);
	full_adder  FA328(carry14[10],sum14[10],P14[10],sum13[11],carry13[10]);
	full_adder  FA329(carry14[9],sum14[9],P14[9],sum13[10],carry13[9]);
	full_adder  FA330(carry14[8],sum14[8],P14[8],sum13[9],carry13[8]);
	full_adder  FA331(carry14[7],sum14[7],P14[7],sum13[8],carry13[7]);
	full_adder  FA332(carry14[6],sum14[6],P14[6],sum13[7],carry13[6]);
	full_adder  FA333(carry14[5],sum14[5],P14[5],sum13[6],carry13[5]);
	full_adder  FA334(carry14[4],sum14[4],P14[4],sum13[5],carry13[4]);
	full_adder  FA335(carry14[3],sum14[3],P14[3],sum13[4],carry13[3]);
	full_adder  FA336(carry14[2],sum14[2],P14[2],sum13[3],carry13[2]);
	full_adder  FA337(carry14[1],sum14[1],P14[1],sum13[2],carry13[1]);
	full_adder  FA338(carry14[0],sum14[0],P14[0],sum13[1],carry13[0]);
	full_adder  FA339(carry15[25],sum15[25],P15[25],sum14[26],carry14[25]);
	full_adder  FA340(carry15[24],sum15[24],P15[24],sum14[25],carry14[24]);
	full_adder  FA341(carry15[23],sum15[23],P15[23],sum14[24],carry14[23]);
	full_adder  FA342(carry15[22],sum15[22],P15[22],sum14[23],carry14[22]);
	full_adder  FA343(carry15[21],sum15[21],P15[21],sum14[22],carry14[21]);
	full_adder  FA344(carry15[20],sum15[20],P15[20],sum14[21],carry14[20]);
	full_adder  FA345(carry15[19],sum15[19],P15[19],sum14[20],carry14[19]);
	full_adder  FA346(carry15[18],sum15[18],P15[18],sum14[19],carry14[18]);
	full_adder  FA347(carry15[17],sum15[17],P15[17],sum14[18],carry14[17]);
	full_adder  FA348(carry15[16],sum15[16],P15[16],sum14[17],carry14[16]);
	full_adder  FA349(carry15[15],sum15[15],P15[15],sum14[16],carry14[15]);
	full_adder  FA350(carry15[14],sum15[14],P15[14],sum14[15],carry14[14]);
	full_adder  FA351(carry15[13],sum15[13],P15[13],sum14[14],carry14[13]);
	full_adder  FA352(carry15[12],sum15[12],P15[12],sum14[13],carry14[12]);
	full_adder  FA353(carry15[11],sum15[11],P15[11],sum14[12],carry14[11]);
	full_adder  FA354(carry15[10],sum15[10],P15[10],sum14[11],carry14[10]);
	full_adder  FA355(carry15[9],sum15[9],P15[9],sum14[10],carry14[9]);
	full_adder  FA356(carry15[8],sum15[8],P15[8],sum14[9],carry14[8]);
	full_adder  FA357(carry15[7],sum15[7],P15[7],sum14[8],carry14[7]);
	full_adder  FA358(carry15[6],sum15[6],P15[6],sum14[7],carry14[6]);
	full_adder  FA359(carry15[5],sum15[5],P15[5],sum14[6],carry14[5]);
	full_adder  FA360(carry15[4],sum15[4],P15[4],sum14[5],carry14[4]);
	full_adder  FA361(carry15[3],sum15[3],P15[3],sum14[4],carry14[3]);
	full_adder  FA362(carry15[2],sum15[2],P15[2],sum14[3],carry14[2]);
	full_adder  FA363(carry15[1],sum15[1],P15[1],sum14[2],carry14[1]);
	full_adder  FA364(carry15[0],sum15[0],P15[0],sum14[1],carry14[0]);
	full_adder  FA365(carry16[25],sum16[25],P16[25],sum15[26],carry15[25]);
	full_adder  FA366(carry16[24],sum16[24],P16[24],sum15[25],carry15[24]);
	full_adder  FA367(carry16[23],sum16[23],P16[23],sum15[24],carry15[23]);
	full_adder  FA368(carry16[22],sum16[22],P16[22],sum15[23],carry15[22]);
	full_adder  FA369(carry16[21],sum16[21],P16[21],sum15[22],carry15[21]);
	full_adder  FA370(carry16[20],sum16[20],P16[20],sum15[21],carry15[20]);
	full_adder  FA371(carry16[19],sum16[19],P16[19],sum15[20],carry15[19]);
	full_adder  FA372(carry16[18],sum16[18],P16[18],sum15[19],carry15[18]);
	full_adder  FA373(carry16[17],sum16[17],P16[17],sum15[18],carry15[17]);
	full_adder  FA374(carry16[16],sum16[16],P16[16],sum15[17],carry15[16]);
	full_adder  FA375(carry16[15],sum16[15],P16[15],sum15[16],carry15[15]);
	full_adder  FA376(carry16[14],sum16[14],P16[14],sum15[15],carry15[14]);
	full_adder  FA377(carry16[13],sum16[13],P16[13],sum15[14],carry15[13]);
	full_adder  FA378(carry16[12],sum16[12],P16[12],sum15[13],carry15[12]);
	full_adder  FA379(carry16[11],sum16[11],P16[11],sum15[12],carry15[11]);
	full_adder  FA380(carry16[10],sum16[10],P16[10],sum15[11],carry15[10]);
	full_adder  FA381(carry16[9],sum16[9],P16[9],sum15[10],carry15[9]);
	full_adder  FA382(carry16[8],sum16[8],P16[8],sum15[9],carry15[8]);
	full_adder  FA383(carry16[7],sum16[7],P16[7],sum15[8],carry15[7]);
	full_adder  FA384(carry16[6],sum16[6],P16[6],sum15[7],carry15[6]);
	full_adder  FA385(carry16[5],sum16[5],P16[5],sum15[6],carry15[5]);
	full_adder  FA386(carry16[4],sum16[4],P16[4],sum15[5],carry15[4]);
	full_adder  FA387(carry16[3],sum16[3],P16[3],sum15[4],carry15[3]);
	full_adder  FA388(carry16[2],sum16[2],P16[2],sum15[3],carry15[2]);
	full_adder  FA389(carry16[1],sum16[1],P16[1],sum15[2],carry15[1]);
	full_adder  FA390(carry16[0],sum16[0],P16[0],sum15[1],carry15[0]);
	full_adder  FA391(carry17[25],sum17[25],P17[25],sum16[26],carry16[25]);
	full_adder  FA392(carry17[24],sum17[24],P17[24],sum16[25],carry16[24]);
	full_adder  FA393(carry17[23],sum17[23],P17[23],sum16[24],carry16[23]);
	full_adder  FA394(carry17[22],sum17[22],P17[22],sum16[23],carry16[22]);
	full_adder  FA395(carry17[21],sum17[21],P17[21],sum16[22],carry16[21]);
	full_adder  FA396(carry17[20],sum17[20],P17[20],sum16[21],carry16[20]);
	full_adder  FA397(carry17[19],sum17[19],P17[19],sum16[20],carry16[19]);
	full_adder  FA398(carry17[18],sum17[18],P17[18],sum16[19],carry16[18]);
	full_adder  FA399(carry17[17],sum17[17],P17[17],sum16[18],carry16[17]);
	full_adder  FA400(carry17[16],sum17[16],P17[16],sum16[17],carry16[16]);
	full_adder  FA401(carry17[15],sum17[15],P17[15],sum16[16],carry16[15]);
	full_adder  FA402(carry17[14],sum17[14],P17[14],sum16[15],carry16[14]);
	full_adder  FA403(carry17[13],sum17[13],P17[13],sum16[14],carry16[13]);
	full_adder  FA404(carry17[12],sum17[12],P17[12],sum16[13],carry16[12]);
	full_adder  FA405(carry17[11],sum17[11],P17[11],sum16[12],carry16[11]);
	full_adder  FA406(carry17[10],sum17[10],P17[10],sum16[11],carry16[10]);
	full_adder  FA407(carry17[9],sum17[9],P17[9],sum16[10],carry16[9]);
	full_adder  FA408(carry17[8],sum17[8],P17[8],sum16[9],carry16[8]);
	full_adder  FA409(carry17[7],sum17[7],P17[7],sum16[8],carry16[7]);
	full_adder  FA410(carry17[6],sum17[6],P17[6],sum16[7],carry16[6]);
	full_adder  FA411(carry17[5],sum17[5],P17[5],sum16[6],carry16[5]);
	full_adder  FA412(carry17[4],sum17[4],P17[4],sum16[5],carry16[4]);
	full_adder  FA413(carry17[3],sum17[3],P17[3],sum16[4],carry16[3]);
	full_adder  FA414(carry17[2],sum17[2],P17[2],sum16[3],carry16[2]);
	full_adder  FA415(carry17[1],sum17[1],P17[1],sum16[2],carry16[1]);
	full_adder  FA416(carry17[0],sum17[0],P17[0],sum16[1],carry16[0]);
	full_adder  FA417(carry18[25],sum18[25],P18[25],sum17[26],carry17[25]);
	full_adder  FA418(carry18[24],sum18[24],P18[24],sum17[25],carry17[24]);
	full_adder  FA419(carry18[23],sum18[23],P18[23],sum17[24],carry17[23]);
	full_adder  FA420(carry18[22],sum18[22],P18[22],sum17[23],carry17[22]);
	full_adder  FA421(carry18[21],sum18[21],P18[21],sum17[22],carry17[21]);
	full_adder  FA422(carry18[20],sum18[20],P18[20],sum17[21],carry17[20]);
	full_adder  FA423(carry18[19],sum18[19],P18[19],sum17[20],carry17[19]);
	full_adder  FA424(carry18[18],sum18[18],P18[18],sum17[19],carry17[18]);
	full_adder  FA425(carry18[17],sum18[17],P18[17],sum17[18],carry17[17]);
	full_adder  FA426(carry18[16],sum18[16],P18[16],sum17[17],carry17[16]);
	full_adder  FA427(carry18[15],sum18[15],P18[15],sum17[16],carry17[15]);
	full_adder  FA428(carry18[14],sum18[14],P18[14],sum17[15],carry17[14]);
	full_adder  FA429(carry18[13],sum18[13],P18[13],sum17[14],carry17[13]);
	full_adder  FA430(carry18[12],sum18[12],P18[12],sum17[13],carry17[12]);
	full_adder  FA431(carry18[11],sum18[11],P18[11],sum17[12],carry17[11]);
	full_adder  FA432(carry18[10],sum18[10],P18[10],sum17[11],carry17[10]);
	full_adder  FA433(carry18[9],sum18[9],P18[9],sum17[10],carry17[9]);
	full_adder  FA434(carry18[8],sum18[8],P18[8],sum17[9],carry17[8]);
	full_adder  FA435(carry18[7],sum18[7],P18[7],sum17[8],carry17[7]);
	full_adder  FA436(carry18[6],sum18[6],P18[6],sum17[7],carry17[6]);
	full_adder  FA437(carry18[5],sum18[5],P18[5],sum17[6],carry17[5]);
	full_adder  FA438(carry18[4],sum18[4],P18[4],sum17[5],carry17[4]);
	full_adder  FA439(carry18[3],sum18[3],P18[3],sum17[4],carry17[3]);
	full_adder  FA440(carry18[2],sum18[2],P18[2],sum17[3],carry17[2]);
	full_adder  FA441(carry18[1],sum18[1],P18[1],sum17[2],carry17[1]);
	full_adder  FA442(carry18[0],sum18[0],P18[0],sum17[1],carry17[0]);
	full_adder  FA443(carry19[25],sum19[25],P19[25],sum18[26],carry18[25]);
	full_adder  FA444(carry19[24],sum19[24],P19[24],sum18[25],carry18[24]);
	full_adder  FA445(carry19[23],sum19[23],P19[23],sum18[24],carry18[23]);
	full_adder  FA446(carry19[22],sum19[22],P19[22],sum18[23],carry18[22]);
	full_adder  FA447(carry19[21],sum19[21],P19[21],sum18[22],carry18[21]);
	full_adder  FA448(carry19[20],sum19[20],P19[20],sum18[21],carry18[20]);
	full_adder  FA449(carry19[19],sum19[19],P19[19],sum18[20],carry18[19]);
	full_adder  FA450(carry19[18],sum19[18],P19[18],sum18[19],carry18[18]);
	full_adder  FA451(carry19[17],sum19[17],P19[17],sum18[18],carry18[17]);
	full_adder  FA452(carry19[16],sum19[16],P19[16],sum18[17],carry18[16]);
	full_adder  FA453(carry19[15],sum19[15],P19[15],sum18[16],carry18[15]);
	full_adder  FA454(carry19[14],sum19[14],P19[14],sum18[15],carry18[14]);
	full_adder  FA455(carry19[13],sum19[13],P19[13],sum18[14],carry18[13]);
	full_adder  FA456(carry19[12],sum19[12],P19[12],sum18[13],carry18[12]);
	full_adder  FA457(carry19[11],sum19[11],P19[11],sum18[12],carry18[11]);
	full_adder  FA458(carry19[10],sum19[10],P19[10],sum18[11],carry18[10]);
	full_adder  FA459(carry19[9],sum19[9],P19[9],sum18[10],carry18[9]);
	full_adder  FA460(carry19[8],sum19[8],P19[8],sum18[9],carry18[8]);
	full_adder  FA461(carry19[7],sum19[7],P19[7],sum18[8],carry18[7]);
	full_adder  FA462(carry19[6],sum19[6],P19[6],sum18[7],carry18[6]);
	full_adder  FA463(carry19[5],sum19[5],P19[5],sum18[6],carry18[5]);
	full_adder  FA464(carry19[4],sum19[4],P19[4],sum18[5],carry18[4]);
	full_adder  FA465(carry19[3],sum19[3],P19[3],sum18[4],carry18[3]);
	full_adder  FA466(carry19[2],sum19[2],P19[2],sum18[3],carry18[2]);
	full_adder  FA467(carry19[1],sum19[1],P19[1],sum18[2],carry18[1]);
	full_adder  FA468(carry19[0],sum19[0],P19[0],sum18[1],carry18[0]);
	full_adder  FA469(carry20[25],sum20[25],P20[25],sum19[26],carry19[25]);
	full_adder  FA470(carry20[24],sum20[24],P20[24],sum19[25],carry19[24]);
	full_adder  FA471(carry20[23],sum20[23],P20[23],sum19[24],carry19[23]);
	full_adder  FA472(carry20[22],sum20[22],P20[22],sum19[23],carry19[22]);
	full_adder  FA473(carry20[21],sum20[21],P20[21],sum19[22],carry19[21]);
	full_adder  FA474(carry20[20],sum20[20],P20[20],sum19[21],carry19[20]);
	full_adder  FA475(carry20[19],sum20[19],P20[19],sum19[20],carry19[19]);
	full_adder  FA476(carry20[18],sum20[18],P20[18],sum19[19],carry19[18]);
	full_adder  FA477(carry20[17],sum20[17],P20[17],sum19[18],carry19[17]);
	full_adder  FA478(carry20[16],sum20[16],P20[16],sum19[17],carry19[16]);
	full_adder  FA479(carry20[15],sum20[15],P20[15],sum19[16],carry19[15]);
	full_adder  FA480(carry20[14],sum20[14],P20[14],sum19[15],carry19[14]);
	full_adder  FA481(carry20[13],sum20[13],P20[13],sum19[14],carry19[13]);
	full_adder  FA482(carry20[12],sum20[12],P20[12],sum19[13],carry19[12]);
	full_adder  FA483(carry20[11],sum20[11],P20[11],sum19[12],carry19[11]);
	full_adder  FA484(carry20[10],sum20[10],P20[10],sum19[11],carry19[10]);
	full_adder  FA485(carry20[9],sum20[9],P20[9],sum19[10],carry19[9]);
	full_adder  FA486(carry20[8],sum20[8],P20[8],sum19[9],carry19[8]);
	full_adder  FA487(carry20[7],sum20[7],P20[7],sum19[8],carry19[7]);
	full_adder  FA488(carry20[6],sum20[6],P20[6],sum19[7],carry19[6]);
	full_adder  FA489(carry20[5],sum20[5],P20[5],sum19[6],carry19[5]);
	full_adder  FA490(carry20[4],sum20[4],P20[4],sum19[5],carry19[4]);
	full_adder  FA491(carry20[3],sum20[3],P20[3],sum19[4],carry19[3]);
	full_adder  FA492(carry20[2],sum20[2],P20[2],sum19[3],carry19[2]);
	full_adder  FA493(carry20[1],sum20[1],P20[1],sum19[2],carry19[1]);
	full_adder  FA494(carry20[0],sum20[0],P20[0],sum19[1],carry19[0]);
	full_adder  FA495(carry21[25],sum21[25],P21[25],sum20[26],carry20[25]);
	full_adder  FA496(carry21[24],sum21[24],P21[24],sum20[25],carry20[24]);
	full_adder  FA497(carry21[23],sum21[23],P21[23],sum20[24],carry20[23]);
	full_adder  FA498(carry21[22],sum21[22],P21[22],sum20[23],carry20[22]);
	full_adder  FA499(carry21[21],sum21[21],P21[21],sum20[22],carry20[21]);
	full_adder  FA500(carry21[20],sum21[20],P21[20],sum20[21],carry20[20]);
	full_adder  FA501(carry21[19],sum21[19],P21[19],sum20[20],carry20[19]);
	full_adder  FA502(carry21[18],sum21[18],P21[18],sum20[19],carry20[18]);
	full_adder  FA503(carry21[17],sum21[17],P21[17],sum20[18],carry20[17]);
	full_adder  FA504(carry21[16],sum21[16],P21[16],sum20[17],carry20[16]);
	full_adder  FA505(carry21[15],sum21[15],P21[15],sum20[16],carry20[15]);
	full_adder  FA506(carry21[14],sum21[14],P21[14],sum20[15],carry20[14]);
	full_adder  FA507(carry21[13],sum21[13],P21[13],sum20[14],carry20[13]);
	full_adder  FA508(carry21[12],sum21[12],P21[12],sum20[13],carry20[12]);
	full_adder  FA509(carry21[11],sum21[11],P21[11],sum20[12],carry20[11]);
	full_adder  FA510(carry21[10],sum21[10],P21[10],sum20[11],carry20[10]);
	full_adder  FA511(carry21[9],sum21[9],P21[9],sum20[10],carry20[9]);
	full_adder  FA512(carry21[8],sum21[8],P21[8],sum20[9],carry20[8]);
	full_adder  FA513(carry21[7],sum21[7],P21[7],sum20[8],carry20[7]);
	full_adder  FA514(carry21[6],sum21[6],P21[6],sum20[7],carry20[6]);
	full_adder  FA515(carry21[5],sum21[5],P21[5],sum20[6],carry20[5]);
	full_adder  FA516(carry21[4],sum21[4],P21[4],sum20[5],carry20[4]);
	full_adder  FA517(carry21[3],sum21[3],P21[3],sum20[4],carry20[3]);
	full_adder  FA518(carry21[2],sum21[2],P21[2],sum20[3],carry20[2]);
	full_adder  FA519(carry21[1],sum21[1],P21[1],sum20[2],carry20[1]);
	full_adder  FA520(carry21[0],sum21[0],P21[0],sum20[1],carry20[0]);
	full_adder  FA521(carry22[25],sum22[25],P22[25],sum21[26],carry21[25]);
	full_adder  FA522(carry22[24],sum22[24],P22[24],sum21[25],carry21[24]);
	full_adder  FA523(carry22[23],sum22[23],P22[23],sum21[24],carry21[23]);
	full_adder  FA524(carry22[22],sum22[22],P22[22],sum21[23],carry21[22]);
	full_adder  FA525(carry22[21],sum22[21],P22[21],sum21[22],carry21[21]);
	full_adder  FA526(carry22[20],sum22[20],P22[20],sum21[21],carry21[20]);
	full_adder  FA527(carry22[19],sum22[19],P22[19],sum21[20],carry21[19]);
	full_adder  FA528(carry22[18],sum22[18],P22[18],sum21[19],carry21[18]);
	full_adder  FA529(carry22[17],sum22[17],P22[17],sum21[18],carry21[17]);
	full_adder  FA530(carry22[16],sum22[16],P22[16],sum21[17],carry21[16]);
	full_adder  FA531(carry22[15],sum22[15],P22[15],sum21[16],carry21[15]);
	full_adder  FA532(carry22[14],sum22[14],P22[14],sum21[15],carry21[14]);
	full_adder  FA533(carry22[13],sum22[13],P22[13],sum21[14],carry21[13]);
	full_adder  FA534(carry22[12],sum22[12],P22[12],sum21[13],carry21[12]);
	full_adder  FA535(carry22[11],sum22[11],P22[11],sum21[12],carry21[11]);
	full_adder  FA536(carry22[10],sum22[10],P22[10],sum21[11],carry21[10]);
	full_adder  FA537(carry22[9],sum22[9],P22[9],sum21[10],carry21[9]);
	full_adder  FA538(carry22[8],sum22[8],P22[8],sum21[9],carry21[8]);
	full_adder  FA539(carry22[7],sum22[7],P22[7],sum21[8],carry21[7]);
	full_adder  FA540(carry22[6],sum22[6],P22[6],sum21[7],carry21[6]);
	full_adder  FA541(carry22[5],sum22[5],P22[5],sum21[6],carry21[5]);
	full_adder  FA542(carry22[4],sum22[4],P22[4],sum21[5],carry21[4]);
	full_adder  FA543(carry22[3],sum22[3],P22[3],sum21[4],carry21[3]);
	full_adder  FA544(carry22[2],sum22[2],P22[2],sum21[3],carry21[2]);
	full_adder  FA545(carry22[1],sum22[1],P22[1],sum21[2],carry21[1]);
	full_adder  FA546(carry22[0],sum22[0],P22[0],sum21[1],carry21[0]);
	full_adder  FA547(carry23[25],sum23[25],P23[25],sum22[26],carry22[25]);
	full_adder  FA548(carry23[24],sum23[24],P23[24],sum22[25],carry22[24]);
	full_adder  FA549(carry23[23],sum23[23],P23[23],sum22[24],carry22[23]);
	full_adder  FA550(carry23[22],sum23[22],P23[22],sum22[23],carry22[22]);
	full_adder  FA551(carry23[21],sum23[21],P23[21],sum22[22],carry22[21]);
	full_adder  FA552(carry23[20],sum23[20],P23[20],sum22[21],carry22[20]);
	full_adder  FA553(carry23[19],sum23[19],P23[19],sum22[20],carry22[19]);
	full_adder  FA554(carry23[18],sum23[18],P23[18],sum22[19],carry22[18]);
	full_adder  FA555(carry23[17],sum23[17],P23[17],sum22[18],carry22[17]);
	full_adder  FA556(carry23[16],sum23[16],P23[16],sum22[17],carry22[16]);
	full_adder  FA557(carry23[15],sum23[15],P23[15],sum22[16],carry22[15]);
	full_adder  FA558(carry23[14],sum23[14],P23[14],sum22[15],carry22[14]);
	full_adder  FA559(carry23[13],sum23[13],P23[13],sum22[14],carry22[13]);
	full_adder  FA560(carry23[12],sum23[12],P23[12],sum22[13],carry22[12]);
	full_adder  FA561(carry23[11],sum23[11],P23[11],sum22[12],carry22[11]);
	full_adder  FA562(carry23[10],sum23[10],P23[10],sum22[11],carry22[10]);
	full_adder  FA563(carry23[9],sum23[9],P23[9],sum22[10],carry22[9]);
	full_adder  FA564(carry23[8],sum23[8],P23[8],sum22[9],carry22[8]);
	full_adder  FA565(carry23[7],sum23[7],P23[7],sum22[8],carry22[7]);
	full_adder  FA566(carry23[6],sum23[6],P23[6],sum22[7],carry22[6]);
	full_adder  FA567(carry23[5],sum23[5],P23[5],sum22[6],carry22[5]);
	full_adder  FA568(carry23[4],sum23[4],P23[4],sum22[5],carry22[4]);
	full_adder  FA569(carry23[3],sum23[3],P23[3],sum22[4],carry22[3]);
	full_adder  FA570(carry23[2],sum23[2],P23[2],sum22[3],carry22[2]);
	full_adder  FA571(carry23[1],sum23[1],P23[1],sum22[2],carry22[1]);
	full_adder  FA572(carry23[0],sum23[0],P23[0],sum22[1],carry22[0]);
	full_adder  FA573(carry24[25],sum24[25],P24[25],sum23[26],carry23[25]);
	full_adder  FA574(carry24[24],sum24[24],P24[24],sum23[25],carry23[24]);
	full_adder  FA575(carry24[23],sum24[23],P24[23],sum23[24],carry23[23]);
	full_adder  FA576(carry24[22],sum24[22],P24[22],sum23[23],carry23[22]);
	full_adder  FA577(carry24[21],sum24[21],P24[21],sum23[22],carry23[21]);
	full_adder  FA578(carry24[20],sum24[20],P24[20],sum23[21],carry23[20]);
	full_adder  FA579(carry24[19],sum24[19],P24[19],sum23[20],carry23[19]);
	full_adder  FA580(carry24[18],sum24[18],P24[18],sum23[19],carry23[18]);
	full_adder  FA581(carry24[17],sum24[17],P24[17],sum23[18],carry23[17]);
	full_adder  FA582(carry24[16],sum24[16],P24[16],sum23[17],carry23[16]);
	full_adder  FA583(carry24[15],sum24[15],P24[15],sum23[16],carry23[15]);
	full_adder  FA584(carry24[14],sum24[14],P24[14],sum23[15],carry23[14]);
	full_adder  FA585(carry24[13],sum24[13],P24[13],sum23[14],carry23[13]);
	full_adder  FA586(carry24[12],sum24[12],P24[12],sum23[13],carry23[12]);
	full_adder  FA587(carry24[11],sum24[11],P24[11],sum23[12],carry23[11]);
	full_adder  FA588(carry24[10],sum24[10],P24[10],sum23[11],carry23[10]);
	full_adder  FA589(carry24[9],sum24[9],P24[9],sum23[10],carry23[9]);
	full_adder  FA590(carry24[8],sum24[8],P24[8],sum23[9],carry23[8]);
	full_adder  FA591(carry24[7],sum24[7],P24[7],sum23[8],carry23[7]);
	full_adder  FA592(carry24[6],sum24[6],P24[6],sum23[7],carry23[6]);
	full_adder  FA593(carry24[5],sum24[5],P24[5],sum23[6],carry23[5]);
	full_adder  FA594(carry24[4],sum24[4],P24[4],sum23[5],carry23[4]);
	full_adder  FA595(carry24[3],sum24[3],P24[3],sum23[4],carry23[3]);
	full_adder  FA596(carry24[2],sum24[2],P24[2],sum23[3],carry23[2]);
	full_adder  FA597(carry24[1],sum24[1],P24[1],sum23[2],carry23[1]);
	full_adder  FA598(carry24[0],sum24[0],P24[0],sum23[1],carry23[0]);
	full_adder  FA599(carry25[25],sum25[25],P25[25],sum24[26],carry24[25]);
	full_adder  FA600(carry25[24],sum25[24],P25[24],sum24[25],carry24[24]);
	full_adder  FA601(carry25[23],sum25[23],P25[23],sum24[24],carry24[23]);
	full_adder  FA602(carry25[22],sum25[22],P25[22],sum24[23],carry24[22]);
	full_adder  FA603(carry25[21],sum25[21],P25[21],sum24[22],carry24[21]);
	full_adder  FA604(carry25[20],sum25[20],P25[20],sum24[21],carry24[20]);
	full_adder  FA605(carry25[19],sum25[19],P25[19],sum24[20],carry24[19]);
	full_adder  FA606(carry25[18],sum25[18],P25[18],sum24[19],carry24[18]);
	full_adder  FA607(carry25[17],sum25[17],P25[17],sum24[18],carry24[17]);
	full_adder  FA608(carry25[16],sum25[16],P25[16],sum24[17],carry24[16]);
	full_adder  FA609(carry25[15],sum25[15],P25[15],sum24[16],carry24[15]);
	full_adder  FA610(carry25[14],sum25[14],P25[14],sum24[15],carry24[14]);
	full_adder  FA611(carry25[13],sum25[13],P25[13],sum24[14],carry24[13]);
	full_adder  FA612(carry25[12],sum25[12],P25[12],sum24[13],carry24[12]);
	full_adder  FA613(carry25[11],sum25[11],P25[11],sum24[12],carry24[11]);
	full_adder  FA614(carry25[10],sum25[10],P25[10],sum24[11],carry24[10]);
	full_adder  FA615(carry25[9],sum25[9],P25[9],sum24[10],carry24[9]);
	full_adder  FA616(carry25[8],sum25[8],P25[8],sum24[9],carry24[8]);
	full_adder  FA617(carry25[7],sum25[7],P25[7],sum24[8],carry24[7]);
	full_adder  FA618(carry25[6],sum25[6],P25[6],sum24[7],carry24[6]);
	full_adder  FA619(carry25[5],sum25[5],P25[5],sum24[6],carry24[5]);
	full_adder  FA620(carry25[4],sum25[4],P25[4],sum24[5],carry24[4]);
	full_adder  FA621(carry25[3],sum25[3],P25[3],sum24[4],carry24[3]);
	full_adder  FA622(carry25[2],sum25[2],P25[2],sum24[3],carry24[2]);
	full_adder  FA623(carry25[1],sum25[1],P25[1],sum24[2],carry24[1]);
	full_adder  FA624(carry25[0],sum25[0],P25[0],sum24[1],carry24[0]);
	full_adder  FA625(carry26[25],sum26[25],P26[25],sum25[26],carry25[25]);
	full_adder  FA626(carry26[24],sum26[24],P26[24],sum25[25],carry25[24]);
	full_adder  FA627(carry26[23],sum26[23],P26[23],sum25[24],carry25[23]);
	full_adder  FA628(carry26[22],sum26[22],P26[22],sum25[23],carry25[22]);
	full_adder  FA629(carry26[21],sum26[21],P26[21],sum25[22],carry25[21]);
	full_adder  FA630(carry26[20],sum26[20],P26[20],sum25[21],carry25[20]);
	full_adder  FA631(carry26[19],sum26[19],P26[19],sum25[20],carry25[19]);
	full_adder  FA632(carry26[18],sum26[18],P26[18],sum25[19],carry25[18]);
	full_adder  FA633(carry26[17],sum26[17],P26[17],sum25[18],carry25[17]);
	full_adder  FA634(carry26[16],sum26[16],P26[16],sum25[17],carry25[16]);
	full_adder  FA635(carry26[15],sum26[15],P26[15],sum25[16],carry25[15]);
	full_adder  FA636(carry26[14],sum26[14],P26[14],sum25[15],carry25[14]);
	full_adder  FA637(carry26[13],sum26[13],P26[13],sum25[14],carry25[13]);
	full_adder  FA638(carry26[12],sum26[12],P26[12],sum25[13],carry25[12]);
	full_adder  FA639(carry26[11],sum26[11],P26[11],sum25[12],carry25[11]);
	full_adder  FA640(carry26[10],sum26[10],P26[10],sum25[11],carry25[10]);
	full_adder  FA641(carry26[9],sum26[9],P26[9],sum25[10],carry25[9]);
	full_adder  FA642(carry26[8],sum26[8],P26[8],sum25[9],carry25[8]);
	full_adder  FA643(carry26[7],sum26[7],P26[7],sum25[8],carry25[7]);
	full_adder  FA644(carry26[6],sum26[6],P26[6],sum25[7],carry25[6]);
	full_adder  FA645(carry26[5],sum26[5],P26[5],sum25[6],carry25[5]);
	full_adder  FA646(carry26[4],sum26[4],P26[4],sum25[5],carry25[4]);
	full_adder  FA647(carry26[3],sum26[3],P26[3],sum25[4],carry25[3]);
	full_adder  FA648(carry26[2],sum26[2],P26[2],sum25[3],carry25[2]);
	full_adder  FA649(carry26[1],sum26[1],P26[1],sum25[2],carry25[1]);
	full_adder  FA650(carry26[0],sum26[0],P26[0],sum25[1],carry25[0]);

	// Generate lower product bits YBITS 
	buf b1(Z[0], P0[0]);
	assign Z[1] = sum1[0];
	assign Z[2] = sum2[0];
	assign Z[3] = sum3[0];
	assign Z[4] = sum4[0];
	assign Z[5] = sum5[0];
	assign Z[6] = sum6[0];
	assign Z[7] = sum7[0];
	assign Z[8] = sum8[0];
	assign Z[9] = sum9[0];
	assign Z[10] = sum10[0];
	assign Z[11] = sum11[0];
	assign Z[12] = sum12[0];
	assign Z[13] = sum13[0];
	assign Z[14] = sum14[0];
	assign Z[15] = sum15[0];
	assign Z[16] = sum16[0];
	assign Z[17] = sum17[0];
	assign Z[18] = sum18[0];
	assign Z[19] = sum19[0];
	assign Z[20] = sum20[0];
	assign Z[21] = sum21[0];
	assign Z[22] = sum22[0];
	assign Z[23] = sum23[0];
	assign Z[24] = sum24[0];
	assign Z[25] = sum25[0];
	assign Z[26] = sum26[0];

	// Final Carry Propagate Addition
	half_adder CPA1(carry27[0],Z[27],carry26[0],sum26[1]);
	full_adder CPA2(carry27[1],Z[28],carry26[1],carry27[0],sum26[2]);
	full_adder CPA3(carry27[2],Z[29],carry26[2],carry27[1],sum26[3]);
	full_adder CPA4(carry27[3],Z[30],carry26[3],carry27[2],sum26[4]);
	full_adder CPA5(carry27[4],Z[31],carry26[4],carry27[3],sum26[5]);
	full_adder CPA6(carry27[5],Z[32],carry26[5],carry27[4],sum26[6]);
	full_adder CPA7(carry27[6],Z[33],carry26[6],carry27[5],sum26[7]);
	full_adder CPA8(carry27[7],Z[34],carry26[7],carry27[6],sum26[8]);
	full_adder CPA9(carry27[8],Z[35],carry26[8],carry27[7],sum26[9]);
	full_adder CPA10(carry27[9],Z[36],carry26[9],carry27[8],sum26[10]);
	full_adder CPA11(carry27[10],Z[37],carry26[10],carry27[9],sum26[11]);
	full_adder CPA12(carry27[11],Z[38],carry26[11],carry27[10],sum26[12]);
	full_adder CPA13(carry27[12],Z[39],carry26[12],carry27[11],sum26[13]);
	full_adder CPA14(carry27[13],Z[40],carry26[13],carry27[12],sum26[14]);
	full_adder CPA15(carry27[14],Z[41],carry26[14],carry27[13],sum26[15]);
	full_adder CPA16(carry27[15],Z[42],carry26[15],carry27[14],sum26[16]);
	full_adder CPA17(carry27[16],Z[43],carry26[16],carry27[15],sum26[17]);
	full_adder CPA18(carry27[17],Z[44],carry26[17],carry27[16],sum26[18]);
	full_adder CPA19(carry27[18],Z[45],carry26[18],carry27[17],sum26[19]);
	full_adder CPA20(carry27[19],Z[46],carry26[19],carry27[18],sum26[20]);
	full_adder CPA21(carry27[20],Z[47],carry26[20],carry27[19],sum26[21]);
	full_adder CPA22(carry27[21],Z[48],carry26[21],carry27[20],sum26[22]);
	full_adder CPA23(carry27[22],Z[49],carry26[22],carry27[21],sum26[23]);
	full_adder CPA24(carry27[23],Z[50],carry26[23],carry27[22],sum26[24]);
	full_adder CPA25(carry27[24],Z[51],carry26[24],carry27[23],sum26[25]);
	full_adder CPA26(Z[53],Z[52],carry26[25],carry27[24],sum26[26]);

endmodule
