module div2_tb();

endmodule